module test_module(y, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10);
output wire [1372:0] y;
input wire [6:0] w1;
input wire [18:0] w2;
input wire [9:0] w3;
input wire [5:0] w4;
input wire w5;
input wire [28:0] w6;
input wire [17:0] w7;
input wire [29:0] w8;
input wire [10:0] w9;
input wire [5:0] w10;
wire [26:0] w11;
wire [21:0] w12;
wire [24:0] w13;
wire [16:0] w14;
wire [10:0] w15;
wire [29:0] w16;
wire [3:0] w17;
wire [25:0] w18;
wire [22:0] w19;
wire [26:0] w20;
wire w21;
wire [6:0] w22;
wire [8:0] w23;
wire [3:0] w24;
wire [24:0] w25;
wire [11:0] w26;
wire [1:0] w27;
wire [24:0] w28;
wire [11:0] w29;
wire [2:0] w30;
wire [4:0] w31;
wire [11:0] w32;
wire [24:0] w33;
wire [27:0] w34;
wire [18:0] w35;
wire [28:0] w36;
wire [5:0] w37;
wire [4:0] w38;
wire [3:0] w39;
wire [12:0] w40;
wire [18:0] w41;
wire [11:0] w42;
wire [3:0] w43;
wire [27:0] w44;
wire [10:0] w45;
wire [8:0] w46;
wire [17:0] w47;
wire w48;
wire [10:0] w49;
wire [14:0] w50;
wire [3:0] w51;
wire [22:0] w52;
wire [1:0] w53;
wire [29:0] w54;
wire [15:0] w55;
wire [10:0] w56;
wire [10:0] w57;
wire [27:0] w58;
wire [24:0] w59;
wire [7:0] w60;
wire [14:0] w61;
wire [17:0] w62;
wire [26:0] w63;
wire [27:0] w64;
wire [4:0] w65;
wire [23:0] w66;
wire [9:0] w67;
wire [9:0] w68;
wire [11:0] w69;
wire [11:0] w70;
wire [19:0] w71;
wire [8:0] w72;
wire [1:0] w73;
wire [5:0] w74;
wire [14:0] w75;
wire [10:0] w76;
wire [8:0] w77;
wire [17:0] w78;
wire [2:0] w79;
wire [10:0] w80;
wire [17:0] w81;
wire [2:0] w82;
wire [21:0] w83;
wire [8:0] w84;
wire [8:0] w85;
wire [10:0] w86;
wire [27:0] w87;
wire [20:0] w88;
wire [12:0] w89;
wire [26:0] w90;
wire [4:0] w91;
wire [25:0] w92;
wire [17:0] w93;
wire [20:0] w94;
wire [25:0] w95;
wire [16:0] w96;
wire [20:0] w97;
wire [17:0] w98;
wire [28:0] w99;
wire [22:0] w100;
assign w11 = w78;
assign w12 = $signed((-13'h10));
assign w13 = ({(w4 < (-21'h7)), (w91 * w38), (^w66), (^~w60), ((26'h8) ? w74 : w55), (w25 ? w30 : (-12'h5)), (w100 >> (36'h10)), ((-6'h11) <= (3'h1d)), (w85 ? (-17'he) : (-19'h1d)), {(20'h9), w73, w3, (9'h19), (-10'h1a), w60, w40, (20'hd), (14'h11), (-3'h1), (-17'h14)}, $signed((12'h9)), ((7'h1b) ? (-1'h1) : w3), (+(17'hd)), (+(14'h3)), ((17'h11) ^ (-15'h13)), (-29'h18), (+w67), $signed((23'h9)), {w42, (-2'h12), w100, (13'ha), (5'h1), w34, w59, w78, (26'hd), w32, w21, (-6'h19)}, $signed((-2'h11)), (+w93), w65, $unsigned(w22), ((-13'h4) ~^ w69), {w71, (-27'h1c), (22'h6), (-18'h15), (26'h18), (21'h17), w16, w69, (23'hc)}, ((-6'he) <= w64), w43, (-(-21'h2)), (w61 ? w93 : (-18'he)), w94} | (w41 >>> $signed((1'hb))));
assign w14 = ((~^(&({(-17'h2), w90, w90, w3, w85, (-6'hc), (4'h1c), w58, (-23'h12), w56, w86, w85, (3'h10), (24'hf), w56, (-23'h3), w46, (13'h19), w41, (-2'h7), w77, (-14'h6), w87, w69} > {w16, (-3'h13), w61, (-13'h8), w7, (11'h6), w84, (-27'h3), (24'h1a), (-1'h12), (-21'h8)}))) === {(^w15), (~&w79), w76, ((2'h1a) ? (-5'h16) : (-31'h9)), (-3'h16), (w20 ? w90 : w50), ((11'h3) ? (7'hc) : w24), (&(-7'h14)), (-28'h17), $signed((12'h4))});
assign w15 = w50;
assign w16 = (-2'h1e);
assign w17 = ($signed(({(9'h6), w67, w75, w19, w25, (13'h7), w71, (16'h9), w48, (-6'h4), (27'h17), (3'h11), w65, (24'h15)} != ((~&(-26'h8)) ? (w73 ? w28 : w10) : (4'he)))) >>> $signed({(-24'h1e), w6, (-23'hc), w98, w84, w53, w26, w63, (6'h1b), (-19'h15), w72, (-3'h3), (12'h8), w63, w72, w87, (-12'hd)}));
assign w18 = (-({w27, (4'h1a), w54, (-15'h17), w80, (5'h1), w100, w6, w46, (9'h15), w77, (-35'h6), w93, w100, w33, w99} ^ w6));
assign w19 = (-19'h5);
assign w20 = $unsigned(((+(14'ha)) <= (13'h11)));
assign w21 = (-30'h12);
assign w22 = $unsigned(((+{(9'h12), w60, w88, (-14'h5)}) < $unsigned($signed(((-5'h0) ? w88 : (-6'hf))))));
assign w23 = $unsigned((-32'h17));
assign w24 = {((w2 ^~ w49) & w82), ((w71 ? w71 : (22'h1c)) | ((14'h8) != w38)), (w32 ? ((-28'h11) >= (-23'h1b)) : $signed((27'h1e))), w55, ($unsigned(w87) ? (-24'hf) : (w60 >= w56)), {w35, (-10'hf), (-25'h12), w58, (14'h1e), (10'h9), w63, (4'h15), w54, (-7'he), (-10'h12), (27'h18), (14'hd), w7, (16'hf), w63, w8, (19'h12), w27, (-16'h4), w26, w55, w74, (4'h5), w8, (-6'h16), (11'h1c), w38, (11'h1a)}, (-24'ha), w37, (25'h3), ($unsigned(w70) != (-3'h9)), (~&$unsigned((-10'h19))), {w8, w96, w36, w33, w100, (-6'hf), (-8'hc), w59, w72, (-14'h1d), (-11'h2), w68, w4, w36, w61, w9, (2'h1), (-17'h16), w30, (9'h13), w89, (-19'h9), w97, w60}, (~^(-25'h12)), {w54, (-3'hc), w56, w45, (10'h17), (-17'h19), w85, w61, (13'h1d), w49, w30, w26, (-12'h5), (-18'h13), (-28'h1a), (27'h19), w7, (20'h10), w78, (-15'h1c), (8'h2)}, $unsigned((w98 !== (-10'h1e))), w57, {(-30'ha), (-3'h17), (29'h2), (-26'h13), (-32'h3), (-22'h5), (5'h3), w69, w85, w9, w95, (-19'ha), (-29'h16), w34, (-19'h1e), w77, (-9'h14), w49, (31'h10), w87, (-10'h19), (-4'h3), (6'h4), w39, w4, w56, (-14'h1e), w92}, ({(11'h5), w47, w41, (23'ha), (-15'h0), (-4'hd), (16'h1d), (-9'hb), (18'h3)} ? (-21'h12) : {w67, (-20'h15), w32, w90, w52, w88, w35, (19'h16), (-12'hf), (15'h1a), w42, w75, w36, (-29'h8), (34'h1), w87, (-31'ha), w57, w8, (-27'h9)})};
assign w25 = ((3'h4) ? (({(26'h1b), (10'hf), (-9'h5), (21'h1b), w90, w59} >> {w74, w53, w76, (22'hd), w86}) ? ({w54, w41, w26, w37, (-28'h3), w9, (-11'hd), (-22'h6), (18'h1), (16'h1a), w98, w3, (22'hc), (-19'he), w60} ? (&(-4'h1b)) : (-4'h18)) : (w5 < (-(-6'h10)))) : {{w57, w3, w86, (-6'hc), w99, (9'h18), (23'h2), w3, w26, (-16'h4), w63, (24'h2), w83, (29'h14), (-30'h1d), w71, w96, (5'h16), (17'hd), (7'h14), (-2'h15), (-20'h5), (28'h19), w64}, {(-29'h1e), w30, (-24'h19), (24'hf), (-11'hc), (7'hd), (1'h5), (23'h3), w49, w98, (25'h15), w80, w98, w61, (21'h7), w61, (-28'h15), w61, w93, (22'hd), (-12'hb), (20'h11), (-24'h6), w6, (-13'hd), w65, (31'h1c), w71, w47, (13'h1)}, ((10'h10) > (27'h1)), (~|(-11'h17)), $unsigned((-2'h11)), $signed((-4'h12)), (-29'h7), (-19'h6), (~|w80), w86, (w51 ? w75 : (10'h7)), {(-17'ha), w48, (7'h12), w67, (23'he), (11'h2), w1, w96, w88}, w62, {(23'h1d), w83}, (+w5), ((9'h19) ~^ w76), w51, ((21'h10) + w99), (&w2), (^(-6'h15)), (-w56), ((20'h5) ? w64 : w63), w50, (w70 ? w95 : w87), w83, (9'h1b), w9, $signed((24'h14)), (+(-20'hd))});
assign w26 = (($signed((-12'h0)) <= w32) && w72);
assign w27 = $signed((^(-15'h1d)));
assign w28 = $signed($signed((8'h1c)));
assign w29 = (^(~|$signed(w9)));
assign w30 = $signed({w3, w79});
assign w31 = $unsigned($signed($signed($signed(w82))));
assign w32 = ((({w7} * $unsigned($signed(w62))) ? w57 : $unsigned((|(+w1)))) & (-35'h0));
assign w33 = (~|w78);
assign w34 = (30'h17);
assign w35 = ((({w1, w4, (-4'h7), w73, (-26'hb), (-22'h12), w8, (-20'h11), (-24'he), w98} || ($signed(w7) ? (17'h12) : (w74 ? w68 : w100))) ~^ (((w10 << w1) >>> {(-22'h8), w45, (-9'hf), (-28'h1), (-12'hf), (16'h1b), (29'h17), (-19'h6), (3'h10), w94, w10, (-32'h2), (-14'h3), (19'h2), (-19'h1), (12'h7), (-30'h15), w92, (18'h3), w60, w54, w100}) !== (-24'h1))) < w37);
assign w36 = (-(-((&(~&(-22'h16))) & $unsigned($unsigned(w42)))));
assign w37 = (!((~|{(-18'h4), w42, (-27'h7), w60, (23'h11), (24'ha), (30'he), w90, w64, w40}) <<< (-27'h5)));
assign w38 = (24'h13);
assign w39 = (^~$unsigned($signed(w8)));
assign w40 = {$unsigned((w83 ? (-6'h1d) : (26'h14))), (~|(w58 ? w98 : (-15'h1e))), (w81 * $signed(w43)), (3'h3), (w60 ? $signed((-6'h10)) : ((28'h18) ? w47 : (-20'h5))), (-14'h15), ((~^(15'h3)) ? (10'h5) : (-2'hf)), $signed(w10), w9, (16'h16), (((-32'ha) ? w83 : w72) ? (+(32'h1)) : (^~(2'h7))), ((19'h13) ? w76 : (-3'h12)), (-20'h13), ($unsigned(w89) ? (-19'h18) : (12'h11)), $unsigned({(-31'h0), (1'h1d), w67, w88, w56, (11'h14), w59, (-23'h5), (-30'h8), (4'h6), w81, (-29'ha), (5'hc), w54, w99, (-3'h3), (-14'h5), w49, (16'hd), (22'h1), w45, (-28'h6), w2, w83, w45, (30'h1d), w87}), (^~(6'h5))};
assign w41 = w5;
assign w42 = {w88, ((w57 << (14'h1)) >= $signed(w8)), w72, $signed((-30'h6)), ($signed(w90) >>> w74), ((-1'h12) ? ((9'h4) ? w73 : (24'hd)) : (-17'h14)), {(-17'h7), w52, w100, w87, w43, (23'hd), (2'h17), (19'h16), (-10'h16), (17'h7), (-24'hb), w75, (5'h5), w68, w53, (-13'h17), (-15'h0)}, w52, ({(13'h4), (18'h10), w50, (5'h16), (-28'h10)} ? (-25'h6) : $signed((12'hf)))};
assign w43 = (($unsigned(w90) ? ((w89 ? (23'h18) : w44) ? ((-2'h3) >= (20'h1c)) : $signed((13'h1e))) : ({w61, (-23'h10), w57} ? (w51 >= w2) : w53)) ? $signed({w65, (1'h19), w98, w70, (9'h1d), w76, w88, w70, w51, (27'h3), w71, (-5'h2), (12'h10), (24'hb), w48, w72, w8, (-10'h1c), (-11'hf), (-15'h3), (-5'h1d), (19'hd), (6'h3), (-15'h1b), w94, w63, w1, (-10'h19), (-17'h15)}) : (+{(-9'hb), (10'hf), w94, (14'h1b), (19'h1b), (-2'h1), (16'h17), (-30'h2), w94, w69, w91, (-10'h3), w89, (-7'h9), (-30'h1), (12'h17), (-6'hb), w84, w79, w97, w70, (19'h5)}));
assign w44 = ((w48 ? $signed((17'h14)) : {(13'h6), (-18'h18), (23'ha), (3'h1b), (10'he), w65, (10'h1d), (30'h2), w45, (-23'h1e), w53, w57, w65, (27'h8), (14'h18)}) ? {(-2'h7), (w61 !== w2), (!w68), (^(16'h18)), (~|(14'h3)), (30'h16), w59, {w100, w94, (-25'h1a), (8'ha), w3, (-18'h5), w84, (-25'h0), (-17'h3), (20'h1), w8, (21'hd), (21'h18), (30'h1e)}, (w82 < (16'hc)), (-19'h0), (w93 == w10), ((-2'h17) ? w7 : w7), (17'h1), ((30'h2) ? w53 : (24'he)), (w52 * (30'h14)), (26'h13), {(11'h9), (7'h16), w75, w3, (1'h5), (30'hf), (-24'hd), w79, (23'h18), (-18'hf), w1, w52, w74}, (11'h1c), $unsigned((-30'h2)), (^~(-12'h18)), {(-22'h1b), w51, w81, (-7'h1c), (-19'h19), (18'h17), w78, (-13'h11), w97, (-24'h1a), (-22'hf), (-13'h18), w7, (-25'hd), (-31'h13), (5'h5), w100, w5, w76, (-3'h1c), w75, (25'h6), (12'h19), (13'h8), (12'h8), (10'h6), w77, w84}, (^w72), (9'h7)} : {(w68 ? (7'hf) : (2'h1b)), ((-3'h17) <= (31'h10)), (w8 | (-19'h2)), (w50 ^~ (-29'h9)), (w69 ? w95 : w97), w62, w98, (-11'hb)});
assign w45 = (-12'h6);
assign w46 = $unsigned((-4'h0));
assign w47 = (w87 ? (-12'h6) : {((13'h2) & w48), $unsigned((27'h11)), w74, (w56 == w55), (~^(4'h1e)), (-27'h1), (w50 ? w5 : (19'h3)), (w91 === (-26'hc)), $signed(w78), ((25'he) <<< w75), {w81, w58, w76, (-24'hf), w2, w65, (36'h3), w78, (15'h9), (18'ha), w64, w84, (-5'h1d), w60, w52, (29'hf), w53, (-24'h16), w48}, (3'h11)});
assign w48 = w100;
assign w49 = $signed({((18'h14) ? (32'hf) : (-3'hf)), (-14'hd), {w66, w95, w79, w71}, w98, w53, (^w3), {w80, (-15'h0)}, $signed(w73), $signed((-16'h1d)), ((-31'h1c) && w89)});
assign w50 = {(((-5'h5) | (-17'h3)) ? (+w57) : w65), $signed((16'h1d)), (20'h4), (-w75), $unsigned((-24'h15)), w73, $signed({w52, w65, w69, (16'h6), (28'h9), (-5'hb), w10, (-15'hf), (14'h1c), (-15'he), (-16'h13), w4, (-26'h17), w89, (31'h15), w10, (-31'h1d), (11'h18), (28'h1a), w68, (15'hd), w2, (-10'h12), (-10'h14)}), {w61, w85, (-22'h10), (24'h3)}, w86, {w10, (9'h18), (13'h6), w6, w98, (-1'hc), w63, (9'h1e), w84, (14'h12), (-26'hf), w60, w94, (-20'h17), w88, (-23'h1d), (-12'h1c), w60, (24'h10), (2'ha), (-1'h12), (-8'h16), (-32'h15), w59, w55}, (-13'h14), (~|w1), {(-30'h14), (-24'h1c), w81, w81, (-17'h7), w56, w87, (-32'h1b), w98, w87, (24'h1), w9, (27'h13), w90, (-19'hf), (6'h18), (8'h6), w6, (-28'h1e), (26'h1), (29'h11), w71, (6'h1b), (-13'h3), (8'h18), (-3'h1a), (20'h3), (6'h7), (-19'h1b), w79}, w95, (12'h4), $signed((w3 & w7)), (~&$signed((8'h16))), (-12'h8), (-3'h1a), (|(w51 >= w100)), w69, w69, ({w76} ? w89 : w51), (|((-4'h13) ? (-2'h1b) : w61)), (-3'h18), (w91 ? {w67, (-27'h1e), w73, (-25'hd), w95, w56, w62, w55, (31'h14), w87, w90, (11'ha), w80, (-19'h16), (25'h2), w67, (14'h3), (14'h1b)} : $unsigned((1'h9))), ($unsigned(w6) >> (w7 > w94))};
assign w51 = $signed({{w5, (21'h1e), w3, (14'h1b), w97, w69, w5, w68, (30'h14), w71, (-10'hd), (-17'h1c), w57, (-17'h14), w73, w86, w57, (12'hd), w74, w99}, (-11'h0), ((-9'h1a) ? w3 : w72), (w100 << (20'h1)), $unsigned((12'h17)), (15'h2), (4'he), (~^w10), ((11'h1c) > (-22'h1)), {(-13'hc), (-26'h7), (-19'hb), w97, w75, w95, (8'h1), (-12'h13), (-20'h12), w8, (33'hc), w5, (-27'h10), w8, (8'hd), w67, (-1'ha), (-9'h17), w57, (29'h19), w88, (22'hc), (-6'h12), (-9'he), w67, w52, w87}, ((1'h1a) ? (3'h1a) : (14'h18)), ((-8'h1e) ? (-5'hb) : (-5'h14)), (-25'h17)});
assign w52 = w86;
assign w53 = {(~&{(-17'h18)}), ($unsigned((-28'h14)) != w9), $unsigned(((8'h4) ? (21'h18) : w79)), {w97, w91, (27'h1), w92, w61, (-9'h5), w6, w84, w54, (27'h1c), w96, (9'h1a), (22'h1a), w75, w62, w55, (-4'h3)}, $signed(((7'h13) ? (19'hf) : (22'h4))), ((26'h6) ? ((14'h14) <<< w85) : {w4, w10, w76, (-28'h9), (-28'h8), (20'h1b), (-12'h15), w78, w5, (14'h10), (-27'h14), w64}), {w8, w94, w74, (-28'hc), w99, (-23'h18), w74, w84, w100, (16'h6), (17'hb), w69, (-28'h4), (-30'h8), (-8'h17), w88}, (((16'h7) ? w5 : w74) ? (~&(19'h16)) : {(-6'h7), w77, (21'h1a), (-26'h7), (-10'hd), w4, w73, (14'h1)}), (w77 ? {w1, w85, (-15'h1a), (-29'h2), (-20'h2), w72, w2, w73, w79, (9'hd), (-31'h13), (20'h15), (-13'h14), w91, w80, w9, (8'h15)} : (~&(10'ha))), (2'h16), {w57, w89, (-4'h5), (28'h11), (-9'h6), w67, w83, w64, (-10'h19), w56, (20'h8), w6, w91, (-14'hc), (6'h6), (-6'h0), (-9'h1), w70, (-4'h16), (33'h1a)}, $signed((-33'h1)), (8'h2)};
assign w54 = ((((((21'ha) >> w58) == ((-17'he) ? w92 : w91)) ? {w72, w86, w60, w96, (11'h15), w76, (4'h9), (-23'h1), w74, w78, (26'h17), w100, w100, (12'h15), (-7'h4), w4, w88, w74, w95, (1'h18), w9} : $unsigned((w100 ? w70 : w63))) ^~ w95) | {((10'h1d) + w62), $signed((15'h1a)), (w71 ? w55 : (23'h13))});
assign w55 = $signed((1'h4));
assign w56 = ($unsigned({(-28'h1), (8'h1b)}) ? (|(28'h1b)) : (-1'hb));
assign w57 = ((w82 ^~ $unsigned(w66)) || (^~$unsigned((-23'h1d))));
assign w58 = w6;
assign w59 = (~^(27'h14));
assign w60 = w74;
assign w61 = ($unsigned(((&(-24'h6)) ? ($signed(w76) < (1'h4)) : ((w90 ? w81 : w4) || w65))) <<< ((({w80, (2'h15), (-31'hd), (-8'h17), (17'hc), w81, (26'hb), w95, w78, w97, w88, (24'h17), (9'h1d)} > $unsigned((-8'h1))) || (((-7'h13) ? (-30'hd) : (-7'h17)) ? ((14'h1e) === (23'h1c)) : (w89 ? w9 : w76))) == (17'h13)));
assign w62 = (8'h1b);
assign w63 = {w76, ({(-14'h2), w88, (31'h1), (19'h3), (-16'h2), w1, w3, w9, w99, w83, (25'hb), w97, (-20'h9), w95, (8'h18), w99, w88, (-11'h8), (-26'h18), (-18'hf), w70, w92, w80, (-26'hd), (28'h6), (-15'hf), w89, (4'h8), (-1'hb), w6} ? $unsigned(w78) : $unsigned(w67)), (-12'hf), w99, (-1'h11), ((w9 ? w2 : (15'h12)) ? {w9, w7} : {(11'h4), w10}), ((-25'h1e) >>> (w73 !== (-26'h4))), (-16'hf), (^{w92, (32'h19), (-23'h1), w4, (-15'h6), w86, (-27'h19), (20'h19), (26'h16), (7'ha), (11'h18), (-27'h1), w91, (22'h11), (-18'h4), w89, w81, (-17'h1e), w80, w69, (-7'h9), w82, w88, (-6'h16), w92, (21'h8), w73, (-20'h6), w81, (8'hd)}), (7'hb), ((w65 ? (22'hf) : (-15'h10)) ? (w91 ? (-15'h9) : w4) : w77), ((-25'he) ? (-2'h13) : (w5 ? w7 : (-7'h15))), (~|((-14'he) ? (-2'h4) : w75)), w91, ($unsigned((-14'hb)) == (w66 ? (-9'h1b) : w77))};
assign w64 = (3'h14);
assign w65 = {(29'h10), (((30'h6) ^~ w87) != ((25'h3) <<< w94)), (-29'h6), $unsigned(((-1'h4) <= w73)), w97, $unsigned(w92), $signed(w76), ({w3, (15'h17)} ? ((-24'h8) ~^ w83) : (~|w76)), w97, ((-31'h1b) ? ((14'h3) ? (26'h1e) : (-28'h9)) : w86), ((10'h7) <<< (~|w75))};
assign w66 = {(+((23'hc) + (16'h10))), $unsigned((w94 | (13'h9))), (-19'h8), {w97, w7}, w98, w89, $unsigned((-w73)), ((~^w9) ? w10 : (w75 & w81)), {(-29'h1d), (18'h3), (-16'hc), w9, (25'h7), (-9'hd), (25'h10), w86, w100, (-24'hc), (-1'h13), w9, (-16'h14), w6, (-30'hb), (31'h10), w100}, (~&$unsigned(w99)), ((~^w1) ^~ $unsigned((8'hc))), (~^(w96 >> w6)), (-7'h18), $unsigned({(10'hb), (-6'h10), (-20'h17), w10, (17'h10), w70, w81, (18'h7), (-23'h9), w100, w88, (11'hc), (-9'h7), w72, (-6'h16), (-25'h3), (-13'h12), w99, w4, (-8'h12), w86, (10'h1e), (13'h6), w67, w4})};
assign w67 = $signed({w90, $unsigned(w69), (w8 < w88), (18'h4), w83, (w93 !== w88), (&w91), (!(25'h9)), (-16'h9), {(12'h5), w99, (-5'h19), w96, w92, (-20'hf), w81, w72}, (21'he), w91, w5, ((11'h2) ? w75 : (-12'hd)), {(17'h9), (9'h2), w96, (-25'h9), (-7'h9), w87, (28'hc), w5, (-12'h4), (-19'h1c)}, (w87 ^~ w79), (w5 !== w86), ((19'h12) >= w77), $signed((27'h19)), ((23'h12) >= w90), (w80 ? (26'h1d) : (21'h3)), w94, (-23'h3), w2, w93, {w8, (7'h1), (-12'h1b)}});
assign w68 = (^~$unsigned(w96));
assign w69 = (+(+w6));
assign w70 = (~|w10);
assign w71 = (4'he);
assign w72 = (((~&((-25'h15) || w97)) ? ((-22'h5) ? (-4'h3) : (^w7)) : w100) ? (-24'h1d) : (-24'he));
assign w73 = w6;
assign w74 = (2'h10);
assign w75 = ((~|{w98, w3, (-19'h8), w95, (30'h1c), w7, w92, (7'h6), (-27'hb), w99, w82, w91, (-9'h18), (25'h18), w90, w82}) <<< w9);
assign w76 = w8;
assign w77 = {{(17'h8), (-9'h0), (-17'h1)}, $signed({(-16'hd), w84, w82, w88, w78, (-23'h2), (28'h1b), (-24'h3)}), ((|w98) == {w6, (-31'h1b), (17'hd), w95, w7, (-15'h1a), w89}), {w4, (-18'h1d), w98, w95, (2'he), w99}, (-(!w100)), w82, ((30'h1e) | (^w3)), w5, $signed({(31'h1e), (13'h9), w81, (29'h10), w79, w82, w5, (-11'h16), w84, w80, (-10'h12), (8'h8), (-29'h8), w98, (-5'h17), w99, w92, w90, (-13'h1), (-20'h9), (-24'h1c), w82, w97, w89, w88, w81}), {w94, w78, w83, w92, (24'hc), (5'h19), (8'h1c), w87, w90, w91, w81, (20'hd), w6}, (17'ha), (1'h1a), {(-5'h1), w5, (21'h19), w86, (-16'he), w79, w93, w7, w94, w95, w83, w79}, (!{w78, w8, (-12'h7), (7'h2), w92, (-25'hf), (-30'h8), w7, w86, (26'h8), w93, (-1'h11), w98, w95, (-14'h0), w1, (25'he), (-12'hd), (-12'hf), (-13'h1d), w85, w84, w82, w86, (-29'h15)}), {(-30'ha), w79, w78, (-16'h10), w94, w86, w92, w1, (12'h19), w7, (11'h1d)}, {(-19'h1), w82, (2'h17), w7, w89, w80, (19'hf), w81, (23'h1b), (6'h9), (10'h1e), (15'h4), w79, (-34'he)}, (-14'h1c), (-18'he), (~&$signed((5'he))), (30'h1c), w87, ({w100, (-13'h1a), w96, (18'h1b), (14'h14), w88, (29'h15), (26'h14), (4'h19), w99, w92, (-15'h10)} || (w86 ? w91 : (-26'h4))), {(20'h11), (-9'h17), (1'h15), (15'h1c), (-15'hd), (24'h10), (10'hd), (-11'h12), w99, (23'h19), w4, (-6'h9), w8, (15'h1a), w79, w100, w88, (-27'h1b)}};
assign w78 = (~|({(-22'h19), (5'h7), w99, (-27'h5), w93, w100, w88, (-10'he)} ? (17'h6) : ((11'h19) ? ((23'h5) ? (6'hf) : w86) : (~&(-3'hf)))));
assign w79 = (+(29'h15));
assign w80 = {$unsigned(w7), w86};
assign w81 = $signed((+(-31'h16)));
assign w82 = (&(w6 ? w98 : ((-7'h4) <= (~^$unsigned((30'h16))))));
assign w83 = (+(|(((-32'h10) << ((-16'h18) * w94)) ? (w87 ? w7 : w8) : (w92 <<< ((-29'h12) ? (-3'h1d) : (3'h2))))));
assign w84 = {{(-19'h18), w10, w8, (6'h2)}, w94, (18'h5), (!((17'h1c) ? (-18'h6) : (4'h1))), {(-18'h8), (12'hf), (-2'h19), (-25'h14), w9, (18'he), (-3'h9), w99, (27'h19), w99, (23'h13)}};
assign w85 = $unsigned({(-22'h1d), (^w100), {w95, (-7'h4), (13'h13), w1}, {(-29'h16), w94, (-4'h5), w89, (23'h10), (-20'h4), (3'h7), w6, (4'hb), w95, (-5'h11), (-7'h5), w8, (-23'hb), w4, w90, (25'ha), w8}, w2, {w94, (17'h15), w93, (-3'h7), w93, (30'h19), w99, w3, w8, w4, w96, (11'h4), w1, w94, w95, w92, (16'he), (7'h1a), (16'h14), w87, (12'h8), w92, w7, (-5'h1b), (-27'hf), (28'h11), (-31'h7), w6, w96, (19'h16)}, {w2, (-6'h4), (3'h1a), w92, w87, w91, w8, (-17'h15), (-23'h9), (18'h8), w92, w89, w10, (16'h12), (21'h19), (-16'h14), (1'h1c), (-11'he), w4, w1, w90, (26'h4), (5'h10), (-10'h15), w89, (-10'h1), (9'hf), w87}, ((21'h11) === (-9'h18)), $unsigned((-21'h13)), (22'h17), (w94 ? w6 : w93), (w9 ? w94 : w92), $signed(w10), (&(-28'h18)), ((-12'h0) ~^ (-5'h16)), (22'hd), (-16'h1e), (-6'h3), w3, {w87, (-24'h1a), (22'h8), w9, w10, (-18'h10), (-2'ha), w1, w100, w6, (-3'h1b), w3, (-15'h14), (23'h1d), w4, (-7'h6), w87, w10, (-19'h16), (12'h1c), w4, w95, (12'hc), w3, w1, w3, (-7'he), w9}, $signed((17'h3)), $signed((-16'hb)), (~&w8), (w87 ? (-23'h19) : w7), {w91, w88, w87, (-15'h0), (27'h13), (-28'h0), w94, (-1'h5), w95, w5, (-24'h10), (-6'hd), w94, (7'h14), (-21'hf), w91, w97, (-30'h3), w97, w96, w7, w93, (-26'h11)}});
assign w86 = (-$unsigned(($signed(w2) >= ((w3 !== w96) ~^ ((-30'h5) & w88)))));
assign w87 = {{(13'h16), (23'h1b), w90, (-5'h17), (30'h16), (11'hc), w94, (-20'h17), (-8'h1b), w3, (29'hc), w7, w90, (-1'h1a), (28'h7)}, w6, $unsigned((14'h1c)), ((~^(-13'hc)) ? (~|(2'h7)) : (^~(2'h1b))), {w94, (-16'h14), (25'he), w91, w10, (19'hd), (8'h18), w96, w10, (-28'he), (-16'h11), (23'h15), (14'h1c), w100, w3, (-18'h14), w90, (-3'h1d)}, (^((-3'h19) > (-12'hf))), w95, {w2, (19'h2)}, $signed((-(33'h9))), w97, (+(^~w93)), (|((-28'h0) ? w3 : w92)), $unsigned((&(-2'h1c))), $signed(w4), w100};
assign w88 = {{(-19'h9), w96, (22'h3), w94, w99, w91, (-10'h12), (-7'h1b), (6'h17), (9'h1c), w100, w90, (-25'hf), (13'h13), w5, w6, w90, w91, (-14'h19), (-29'h1e), w98}, (w4 != (18'h1e)), ((w3 ^ w97) < (!(17'h1))), {w92, (-9'h15), (-24'h15), w10, w91, w99, w99}, {w91, (-28'h8)}, {(17'h8), (25'h13), (31'hc), (27'h18), w1, w2, (8'h1), (16'hd), (-25'h4), (13'h1a)}, {(1'hf), (28'h15), (-25'h7), (7'h14), (4'h1b), (-23'h14), (4'h8), (4'h7), (27'h4), w95, w97, w1, (31'h10), (23'h1), w90, w91}, ((20'h9) <= w10), $signed($unsigned(w1)), $unsigned(w90), {(-13'h17), (24'h15), (-23'h13), (-1'h2), w99, (-29'h11), (-18'h1d), (29'h16), (16'h11), (-4'h2), (-29'h3), (27'h1b), (12'h1b), w97, (-28'h13), w95, (3'h3), (14'h12), (-10'h1a), w1, (1'h7)}, (((8'h1e) ? (29'h3) : (25'h4)) <= (-30'h5)), (!((-30'h1b) ? (10'h1c) : w2)), ((w91 == (15'he)) ? (^(1'h7)) : (w96 < (-15'h16))), ((w4 ? w89 : (-29'ha)) ? (~|w95) : {(-28'h16), w1, w93, w92, (30'h1e), (-21'h1d), w6, (25'h1e), (16'h18), w8, w96, w98, w99, (-30'h1c), (-6'h2), w4, (-22'h6), (-18'h3), w10, (-18'h1a), w89, (25'h8), (-17'hb), w2, w98, w94}), ({(7'he), (28'h17), w92} ? {w91, w97, (9'h8), (24'he), (-30'hf), (-4'h12), w2, w2, w90, (7'h1), w7, w9, w6} : w94), $unsigned(((8'hb) ? w4 : w6))};
assign w89 = ($signed((^w94)) ? ($signed((12'he)) ? (-29'hd) : (-28'h16)) : (~^(-21'h13)));
assign w90 = (({(29'h9), w93, w98, (9'h2), w6} ? (10'hd) : (17'h1)) ? $unsigned(((-30'h1d) || (~|w96))) : ({w7, (2'h9), (5'h1e), w97, (-26'h16), (24'h14)} >= (17'h5)));
assign w91 = ((27'h1d) > ($signed(((7'h10) !== (-30'h19))) ~^ {w92, (-30'h1d), (-12'hd), (30'he), (-7'hc), (-25'h16), w93, (-20'h1a), w1, w1, (-1'hc), (-28'h1c), w92}));
assign w92 = ({{w1, w99}, (&(-6'hb)), (-19'hd), (w93 && (-11'hb)), (w94 ? w97 : (-2'h9)), ((-30'h8) ? (-8'he) : (-24'h2)), {w94, (-19'h17), (7'hf), w97, (5'ha), w9, w10, w93, w2, (-28'h0), (-19'hb), w93, w93, w93, (20'h11), (24'h5), w3, (-1'h15), (-4'h17), (27'h13), w96, w7, w95, w94, w93}, (^(-20'h10)), ((-3'h16) > w100)} ? (($unsigned((-30'h1b)) <<< (6'h19)) ? ((~^(23'ha)) == (w98 ^ (-10'h1))) : (20'h16)) : {((28'h4) != w8), (~^(18'h9)), $signed(w97), w1, w94, $signed(w4), w1, ((20'h13) ? (6'h1b) : w97), (^w4), $signed(w97), {(-9'ha), (25'h11), w98, w99, (-19'h18), (12'h1e), (29'h1a), w93, w96, (6'h1), (9'h17), w98, (-13'ha), (-3'h1e), w97, w100, w96, (-21'he), w94, w8}, {(28'ha), (11'hd), (-20'h16), (-13'h3), w98, (-16'h19), w99, w9, w5}, (-29'h13), {w5, (20'ha), w5, w94, (-1'h12), (-26'h12), (2'hd), w8, w6, w94, (-28'hb), (-11'hf), (-7'h2), (27'h16), w8, w95, w2, w8, (1'h10), (-9'h12), (-1'h0)}, ((-20'h5) & w94), {(-30'h16), (-23'h17), w97, (18'h16), (-2'h0), w10, w10, w5, w6, (28'h13), (-19'h0)}, w98, $signed((18'h3)), w8, $unsigned(w97), ((-25'h16) ^~ (-18'h7)), (-15'ha)});
assign w93 = {((+(28'ha)) >>> w2), (-11'h15), $signed(w4), ((12'h7) < w6), (2'h19), (!(-(-30'h19))), ((~&(-15'hf)) ? (^~(12'h17)) : $signed((-4'h1d))), ((^w95) ? $signed(w1) : $unsigned(w5)), $signed((w96 ? (-31'h3) : w100)), w99, w95, w7, (-2'hb), (+w5), ({(-30'h0), w96, w10, (-23'h0), w98, w2, w1, w96, (19'h8), (-22'h18), (3'h1b), (6'h6), w7, w99, (18'h19), (10'he), (16'hf)} ? ((19'h12) ? (-2'h8) : (23'h6)) : $unsigned(w9))};
assign w94 = ((10'hc) ? (~&{w100, w100, (17'he), (10'h1b), (4'h1a), (2'h15), (-4'h4), w3, w1, (-9'hf), (19'h1c), w99, (29'h2)}) : w2);
assign w95 = w3;
assign w96 = $unsigned((-1'h17));
assign w97 = ({(w9 ^ w7), ((-27'he) != w99), ((-19'h17) ? w1 : (23'h1e)), (w10 ? w9 : (1'h11)), (w2 ? (1'hc) : (8'h5)), (-28'h11), (w3 ? w99 : w6), $unsigned(w9), (w98 > (-5'hc)), (-5'h14), ((-20'h0) ^~ (-4'h1b)), {(8'ha), w100, w1, (-3'h1d), w98, w6, w9, (-15'hc), w99, (-18'h4), (-4'h1b), w3, (20'h6), (27'h5), w3}, w99, (~^(-26'h11))} ? $signed(($signed((-7'h1c)) ? (w4 >>> (-2'h4)) : ((-23'h10) && w3))) : {(+(-17'he)), (^(18'h10)), {w2, w98, w7, w98, (-26'h1), w6, w4, (9'hb), (29'h1), (-1'h1e), (-15'h11), (29'h18), (-4'h1a), (23'ha), (24'h14), (17'h10), (28'h14), (32'hc), w99, (-29'hc), (-10'hf), (-24'h11), (31'h19), w2, (-14'h15), w6, w4, (2'hc), w7, (-17'h7)}, (&w100), {(29'h18), (-25'h4), (6'h13), (27'h7), (-22'h18), (-23'h4), w3, (-26'h1), (29'h1d)}, ((19'h1b) ? w3 : w3), (4'ha), $unsigned(w6), ((-19'hc) ? w8 : (29'h9)), w99, (w7 && w4), (|w5), {(7'h4), w1, w3, w98}, w10, ((-2'h13) * w99), (w8 + (-5'h12)), (-17'h16)});
assign w98 = (w4 >> (-11'h3));
assign w99 = w2;
assign w100 = (10'h3);
assign y = {w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100};
endmodule
