module test_module(y, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10);
output wire [1288:0] y;
input wire [17:0] w1;
input wire [11:0] w2;
input wire [24:0] w3;
input wire [2:0] w4;
input wire [26:0] w5;
input wire [22:0] w6;
input wire [2:0] w7;
input wire [10:0] w8;
input wire [23:0] w9;
input wire [5:0] w10;
wire [4:0] w11;
wire [22:0] w12;
wire [7:0] w13;
wire [3:0] w14;
wire [25:0] w15;
wire [11:0] w16;
wire [7:0] w17;
wire [16:0] w18;
wire [10:0] w19;
wire [11:0] w20;
wire [13:0] w21;
wire w22;
wire [22:0] w23;
wire [21:0] w24;
wire [7:0] w25;
wire [10:0] w26;
wire [28:0] w27;
wire [3:0] w28;
wire [25:0] w29;
wire [3:0] w30;
wire [13:0] w31;
wire [23:0] w32;
wire [26:0] w33;
wire [10:0] w34;
wire [11:0] w35;
wire [9:0] w36;
wire [23:0] w37;
wire [14:0] w38;
wire [29:0] w39;
wire [12:0] w40;
wire [24:0] w41;
wire w42;
wire [15:0] w43;
wire [6:0] w44;
wire [5:0] w45;
wire [17:0] w46;
wire [16:0] w47;
wire [3:0] w48;
wire [8:0] w49;
wire [9:0] w50;
wire [14:0] w51;
wire [5:0] w52;
wire [9:0] w53;
wire [2:0] w54;
wire [24:0] w55;
wire [13:0] w56;
wire [12:0] w57;
wire [29:0] w58;
wire [5:0] w59;
wire [10:0] w60;
wire [9:0] w61;
wire [24:0] w62;
wire [15:0] w63;
wire [29:0] w64;
wire [7:0] w65;
wire [15:0] w66;
wire [4:0] w67;
wire [11:0] w68;
wire [12:0] w69;
wire [16:0] w70;
wire [2:0] w71;
wire [3:0] w72;
wire [6:0] w73;
wire [10:0] w74;
wire [26:0] w75;
wire [21:0] w76;
wire [28:0] w77;
wire [23:0] w78;
wire [13:0] w79;
wire [5:0] w80;
wire [28:0] w81;
wire [4:0] w82;
wire [7:0] w83;
wire [29:0] w84;
wire [5:0] w85;
wire [24:0] w86;
wire [3:0] w87;
wire [13:0] w88;
wire [15:0] w89;
wire [13:0] w90;
wire [4:0] w91;
wire [28:0] w92;
wire [7:0] w93;
wire [22:0] w94;
wire [8:0] w95;
wire [6:0] w96;
wire [8:0] w97;
wire [26:0] w98;
wire [9:0] w99;
wire [19:0] w100;
assign w11 = {(w60 ? ((-10'h1b) ~^ (-5'h18)) : (24'h15)), (^(w3 ? (-20'h4) : (-3'hd))), {w2}};
assign w12 = (17'h1e);
assign w13 = {(22'h14), $signed((w1 || w14)), (29'h16), (~&{(-6'hc), (25'hf), w67, w40, (-18'h18), (27'h16), w16, (20'h1), (28'h12), w47, (-16'h15), w9, w34, (-12'h15), (24'h1), (-16'ha), (-26'h7), w53, (14'hd), (18'h10), (-6'h0), (-24'h16), (-18'h17), (-15'h19), w14}), (((-3'h15) & w32) ? w54 : ((23'h1e) ? w91 : (17'h1a)))};
assign w14 = ((($unsigned($signed(w78)) | (-29'h1b)) ? w22 : $signed(((-2'h13) ? w20 : w91))) - {(-19'h1), ((31'hd) >> w66), (w70 ? (-5'h1c) : (-16'h7)), w78});
assign w15 = w81;
assign w16 = {w82, {(25'h15), w96, (-13'hd), (6'hb)}, w50, $signed(w67), $signed({(22'h1d), (-5'h11), w64, w90, w91, w10, w32, w96, w30, (31'h1), (-2'h19), (25'h2), (13'h1b), w5, w70, w35, (-23'ha), w41, (29'h6), w91, w29}), (((-25'h11) ? w20 : w67) > (w21 << (-19'h13))), (&$unsigned((21'ha))), $signed(w69), (-10'h11), ($signed((12'h1c)) ? $signed(w90) : $unsigned((21'h13))), $unsigned(((29'hb) ? (-31'h17) : w51)), ((-16'h19) ? (|(24'hf)) : (~|(-2'h18))), (13'ha), {w93, (15'h1), (-3'h18), w19, w25, w50, (-26'h1b), w26, (11'h18), (32'h1), (13'hc), w45, w57, w52, w18, w17, (-4'h15), (-12'h2), (30'h1a), (5'hf), w7, w1, w71, w36, (-2'h15), (28'h9), (20'h1e), (22'h7)}, $unsigned((|(-6'h6))), ((5'h1c) != (-17'h8)), w96, (~^{(-10'h14), (-8'h19), w34, (27'h10), (8'h17), w21}), (|(w26 ? (22'h1d) : (-11'h5))), $unsigned(((-1'h18) ? w50 : (-2'h8))), ((-15'h1b) === (-29'he)), ((w70 >>> (21'hd)) - $unsigned((-23'h0))), {(22'h13), (-29'hf), w32, w72, w17, w34, (14'he), w79, (22'h6), (24'h10), (17'ha), (-3'h1e), (-19'hd), w21, (11'he), (-13'h1b), (18'h11), w83, w78, w97, (4'h11), (-6'h1b), (17'h8), (-17'h12), w7, w42}, (w53 - w86), (~|w6), {w5, (12'h6), w59, w54, (20'h1), (-8'h12), (11'h4), w100, w95, w96, (-8'h6), w28, (-17'h17), (-6'he), w48, (-29'he), w41, w53, (-21'h1e), (29'h3), (-21'h19), w75, w59, w54, w25}, (~|((-12'h1b) * w93)), {w62, w61, (2'h10), (-2'h0), w63, w58, (-3'h11), w57, (-9'hf), (12'hf), w94, (-10'h3), (2'h1c), (20'h1c), (21'h6), w72, w46, w85, (9'h1d), w1, (13'h3), w31}};
assign w17 = (-26'h3);
assign w18 = w48;
assign w19 = (w92 ? ({(-28'h2), (-29'h18), (13'h4), (22'hf), (21'h16), (-15'he), w89, w88, w77, (-32'h1a), (6'hc), w20, (6'h16), (-8'h17), w45, w78, (-6'h7), (-31'h1a), (-8'he), w93, w59, w92, w32, w8, w50, (-9'h19)} === {(6'h4), w61, w68, w68, (12'h1a), w98, (-26'h1d), (16'h8), (-34'h19), w59, w54, (28'h1a), w98, (4'h9), (4'h16), w49, w54, w46, (17'hf), (28'h5), w1, (-26'h1a), w2, (19'h13), w38}) : w64);
assign w20 = $signed({w21, (!(-17'hb)), $signed((12'h1)), (-w93), w94, (6'he), {(24'h6), w41, w53, (3'h1d), (23'h19), (4'h17), (22'h11), (-30'h11), w81, w70, w7, w27, w94}, $signed((5'h5)), (w3 || (29'h18)), (25'h18), w98, ((21'hc) * w43), $signed((18'h10)), ((6'h1e) || w58), {w87, (-30'h10), (25'h1a), (-15'ha), (24'h18), (23'he), (-2'hd), (14'he), w76, (25'he), w98, w30, (18'hf), (23'h16), w61, w78, w4, w73, (-28'h12), (-30'h1c), (-14'hb), w95, w80, w24, (30'hc), w25, w24, w77, (23'ha)}, ((21'he) | (22'hf)), ((-3'hb) && (10'h18)), $unsigned(w46)});
assign w21 = (2'hd);
assign w22 = {w65, w33, $signed(((-3'hb) + (21'h8))), {w54, (17'h2), w1, w3, w40, (24'h10), w93, (-8'h15)}, {(14'h12), w1, w94, w46, (-28'h18), w70, (-28'hd), (-1'h14)}, {(-11'h1d), (23'h13), (-9'h18), (12'h1), w25, (7'h16), (24'h3), w82, (21'h19), (-4'he), (10'hf), (7'h11), w70}, {(-22'hb), w94, w39, w3, w28, w73, (30'h5), (13'h1c), w89}, (2'h5), w68, (!w3), (((9'h9) ? w89 : w78) ? (w47 ? (-4'h0) : w53) : (-14'h9)), {(17'h1b), (16'h17), w55, (-27'h14), w40, w37, (17'h15), (-3'h11), (21'h1c), w83, w28, (-26'h2), w98, w54, (7'hf), w96, (-15'h5), (2'h5), w43, w29, (8'h2), w75}, w3, $signed(((-19'h14) ? w76 : w78)), (~|((7'h12) ? w89 : w9)), (|w69), $signed($signed(w3)), (|w62), ($signed((15'h12)) < {(16'h6), (-1'ha), (-21'h10), w57, (-2'h15), (-15'hc), w80, w99, w23, (16'h11)}), w4, (((26'h9) ? w51 : w92) && w44), ((w95 != (-16'h10)) ? (w99 * (13'h9)) : {(-9'h19), (29'h1), w35}), ((-10'h14) > w31), ((!(-20'h18)) && ((19'h19) ? (-15'h10) : w62)), w51, {(-14'hb), w28, (24'hf), w7, w26, (-14'h3), (-19'h13), w2, w31}, (w72 ? ((13'h10) >> (4'h8)) : (^~w47)), {(28'h19), w64, (-4'he)}, ((w99 - (19'h15)) < w1)};
assign w23 = ({$signed(w45), {w70, (-21'h18), (7'h14), (17'h3), w41, (2'h8), (-2'h12), w52, w81, w26, w47, w45, w7, (-1'h0), w91, (-13'h12), w36, w76, w6, w2, w60, (20'h6), (-28'h3)}, (26'h8), ((-13'h18) <<< w78), (^(-30'ha))} != ({w61, w33, w68, w36, (14'h1a), (-20'h1a), (22'h17), w4, (-9'he), (6'h10), (-30'h1b), w69, (13'h4), (-3'h5), w9, w84, (-16'h10), (-29'he), (-5'h4), w74, (19'h1b), (-7'h0), (-27'he), w56, w53, w58, (6'h1e), w44} ? {(12'h7), (27'h17), w2, w89, w38, (-24'h1d), w46, w47, (-5'h0), w45, (8'h18), (22'h9), (-11'h16)} : $unsigned((^((7'h8) ? (-18'h15) : w71)))));
assign w24 = {(w62 ? (-14'h5) : (26'ha)), (((-23'h5) ? w37 : (-10'h15)) || $unsigned(w1)), $unsigned({(24'hd), w82, w31, (24'ha), (-27'hf), (-27'h1d), (-23'h18), (-5'h1a), (-14'h1b), w55, (11'h1b), (-29'ha), (-2'h3), w63, w59}), (30'h18), {w28, (3'h18), w56, w99, w36, (2'h11)}, w92, (w53 ? w85 : w7), (((-17'h2) ? (2'h15) : w71) ? (w86 && w7) : (w10 ? (-13'h14) : w98)), (-24'h0), $signed((+w61)), {(-16'h9), w39, (-5'h1a)}, (+(-26'h1c)), (~&w32), (~|(w95 && (-7'h1d))), ((22'h1a) === (w27 ? w85 : (-25'he)))};
assign w25 = {$unsigned((-17'ha)), (((13'he) * (-28'h16)) != w26), (&w29), {w52, w89, w41, w36, (-17'h1d), w10, w92, (1'hc), (9'h19)}, ((^(21'hf)) ~^ ((3'h10) ? w1 : (22'h2))), (~|(-5'h13)), w39, ({(24'h11), w69, (19'h13), (6'h4), w41, w82, (-5'he), w39, w96} || (w77 ? w46 : (11'h2))), {(13'h1e), (8'h1e), w48, (8'h6), w4, (30'h1d)}, w82, (~^{(24'hd), w36, (-29'h4), w92, w61, (25'h1b), w84}), $signed((-2'h8)), $signed({w92, (21'h1b), (-15'h1a), (27'hc), (-7'h13), (-19'hb), w67, w39, (22'h8), (-16'h1), (-30'h16), w79, (27'h9), w55, (-6'h2)}), (~^{w6, (-18'hf), w39, w75, (-26'h0), (17'hd), (-30'he), w87, w8, w42, w80, w62}), ({(17'h5), (29'h1c), (5'h15), w60, w44, w91, (-14'h11), w51, (2'h1d), w6, w61, w5, w76, w27, (-5'h4), (11'h2), (29'h19), (-1'ha), (29'h2), (-24'h1a), w26, w38, (-21'h1d), w68, (-8'h18), w57, w52, w29, (3'h10)} >> (w31 ? (4'h1d) : w32)), (^~(w4 ? (23'h1b) : w77)), ({(-29'he), w79, (-2'h1e), w72, (25'h19), (-16'h5), w68, w53, (-18'h11), w63, w98, w79, (28'he), w79, w90, (25'h8), (9'h16), (13'h5), w65, (-6'hb), (-4'h11), (18'h12), (-8'h1d), (-26'h1e)} ? ((-9'h1) ? (20'h5) : w89) : (!w97)), ((~|(20'h1e)) ? (9'h11) : w96), (4'h2), (-14'h12), ((&(-15'hc)) ? $unsigned((-18'h10)) : (w2 ? w76 : (22'h1))), $unsigned(((-6'h2) ? (-12'h14) : w31))};
assign w26 = ((!w7) ^ $signed(w36));
assign w27 = $signed((-7'h5));
assign w28 = ($unsigned((21'ha)) < (-9'ha));
assign w29 = (-21'h17);
assign w30 = (({w68, (26'h1c), w63, (-18'h17), w55, w61, w42, (-22'h0), (-7'h10), (3'h16), w65, (-22'h12), (-19'hc), w63, w80, (20'h9), w98, (3'h1a), w80, (16'h1e), w70, w56} & (-27'ha)) ? (-28'h1e) : (($unsigned((10'hd)) ? w74 : w99) ^ (^((29'h1c) ? w67 : w10))));
assign w31 = {(-8'hd), $unsigned((w86 ? w77 : (26'hc))), {w67, (-16'h7), w92, w89, (4'h1a), (-7'ha), (29'h7), (-9'h6), w59, (24'h7), w37, w1, w68, (14'hb), (26'h15), (-7'h7)}, (~|((3'h1b) || w96)), (!$signed((-22'h14))), (!(|(-13'h7))), ((~^(-21'h8)) ? (w63 & (24'h2)) : {(-9'he), w52, w86, (-24'h1c), w73, w47, w77, (-10'h18), (5'h10), (10'he), w79, w33, w85, w48, w3, (-21'h5), w60, w36, (-11'h15)}), ((27'h1c) ? $signed(w39) : w66), {(5'hc), w86, w84, w45, w45, w64, w37, w70, w65, (4'hf), (-25'h9)}, {w5, (26'h2)}, ((-5'h18) ? (^~(-1'h12)) : (w38 ? (27'h3) : w51)), w56, {w1, (6'h8), w77, (20'h12), (-14'h6), w100}, (~|((8'h1d) | w99)), w47, w2, {w67, (26'h4), (-3'h3), (8'h7), w48}, w91, w68, (&w8), {(-23'h0), (-7'h0), (-32'hc), w36, w7, (-10'h1d), w92, (-18'h15), (6'h1e), (-29'h1c), w97, w40, (33'hd), w91, w46, (31'hb), w99, (-2'hc), w3, w49, w99, (-7'ha), (-4'he), w80, (12'h1e), w43}, w62, $unsigned({w33, w92, w32, (1'h1c), (-25'h1e), (-16'hf), (15'h13), w74, w44, (18'h13), (24'h16), w10, (24'h8), w33, (7'ha)}), (13'h7), {w10, w64, w10, w70, (10'h1e), (6'h2), (29'h18), w83, w44, w2, w78, w63, (30'h8), w44, w73}};
assign w32 = {({w81, (28'hd), (3'h19), w94, (-6'hf), w33, (1'h19), w54} ? ((-3'h1c) >= (3'h1a)) : (-27'h1)), (~|$unsigned((14'h6))), w60, {(22'hc), w64, (-29'ha), w47, (-12'h1a), (-8'h1e), (14'h11), w39, w34, w1, (-20'h3), w74, (-11'h1a), w82, w95, (17'h10), w70, (-17'h0), (-19'h11), (14'h12), (-11'h1d), w2, (10'ha), w66, (26'h1b), w97}, (^{(15'h5), (5'h17), (-33'h1b), w94, w10, w83, (-13'h1c), w5, (-25'hf)}), (~|(w41 * w6)), w4, $signed($signed(w1)), (^(27'h10)), {w62, (22'h19), (-8'h1c), w62, (19'hc)}, {(-17'h4), w8, (17'h17), w40, w65, (-12'h12), (27'he), (15'h10), w40, (-25'h9), w2, w8, w96, w83, w38, w33, w82, (-4'h17), (18'h4), w57, w72, w2, (17'hd), w88, (-2'h15)}, (-27'h1e), (((3'h2) ? w59 : (12'h15)) ? w88 : (22'h15)), {w65, (-26'h15), (-6'h12), (8'hb), (6'h15), (-7'ha), w46, w84, (13'h4), w93, w51, w63, w89, w85, (3'h1d), w37, w47, w86, (-14'h0), (3'h5), (-31'h4), (13'h12), w43, w43, (-2'h4), (29'h16), w98}, ((~|(-12'h4)) ? (|(7'h11)) : (+(-30'h6))), w39, {(-9'h11), (-17'h1), w33, (22'h19), w39, w53, w59, (5'h19), w57, w8, (-3'h12), w94, (-15'h4), (-7'h8), (11'h7), (9'hf), w83, (31'h6), w4, (5'h1a), (-4'hb), (6'hd), (-2'h1c)}, (~&((6'h1a) >>> w5)), (w83 ? ((-9'ha) == (4'he)) : (w41 ^ w56)), w33, $unsigned((!w89)), (19'h4), (-4'h15), w5, ((w66 ? (-27'h14) : w60) * {(3'h1b), (20'hd), w58, w76, (-5'h3), (27'h6), (15'h18), (11'hb), (-26'h10), w78, (29'h16), w81, w51, (4'h1), w5, (-4'h18), (-11'h12)}), ((+w77) ? ((10'h1b) || (27'h12)) : (^w81)), ((20'hb) * ((17'ha) ? w100 : (-13'h1)))};
assign w33 = ({(!(28'h17)), (18'h1d), ((-13'ha) ? (17'h12) : w76), (!(-13'h1c))} ? {{(8'h19), w4, (-18'hc), (-25'h7), w42, w64, (-15'h15), w81, (-12'h13), w68, (-27'h0), w51, (-16'h1e), w99, w64, w45, w91, w63, (32'h16), (-11'h13), (24'h7), w1, (12'h1)}, (16'h8), (27'ha), (|(6'h12)), {(19'hf), w79, (-3'h15), (-28'h1), w79, (-23'h4), (21'h1d)}, (+(13'h1c)), (+w4)} : {(w77 ? w90 : w44), (w60 + (18'h3)), ((12'h1e) ? w58 : (-12'h5)), w9, ((-26'hf) ^ w70), ((-27'ha) ? w37 : w7), (w55 < w38), ((15'ha) ? w9 : (-21'h16)), {(7'h13), w90, w7, (5'hb), (21'h6), w94, (-5'h6), (24'h18), (-19'hc), (18'h6), w92, (-22'h1c), w86, (16'h13), w71, w57, (-22'h18), (11'he), w2, w6, (20'h16), (29'h9), w100}, (w76 ? (-13'h1d) : (-10'h17)), {(8'h4), w41}, $unsigned(w76), (32'h7), (-12'h7), $signed(w2), (w38 ? (-2'h15) : (6'h17)), w88, ((22'h1e) === (20'h18)), $unsigned(w67), (-19'h1a), (11'h1), w66, w88, ((31'h18) ? w1 : (11'h17)), $unsigned(w96), (!w100), {(-22'h19), (9'h1d), w1, w66, w92, w8, (-27'h16), (11'h11), (12'h1e), (1'hd), w42, w41, (-28'h7), (16'h5), w7, w52}, $unsigned((27'h1d)), ((1'h4) >= w61), $signed((20'he))});
assign w34 = w42;
assign w35 = (&(((w42 ? (19'h1c) : (-31'he)) ? (~|(-2'h9)) : {w72, (-4'hc), w65, w73, w7, (21'hc), w87, w8, (-12'h16), w56, (-5'h4), w78, w42, (-19'ha), w8, w63, w5, w51, (-24'ha), (20'ha), (-18'h12), w70, w93, (10'hb), w7, w9, w97, (16'h4), (-15'h1), w36}) ? {(-25'h0), (-2'hf), w54, w89, (-25'h8), w68, (-31'h19), w52, (-19'h10), (-15'hf), (-17'h10), (23'h9), (-19'h13), w48, w37, w80, (-12'h4), w95, (-27'hb), (-24'h12), w71, w36, w52, w42, w48, (7'h10), (-2'h14)} : (8'h7)));
assign w36 = w94;
assign w37 = ((((w73 ? (-22'h12) : w47) ^ ((22'h7) ? w89 : w50)) * ((w88 ? (10'h6) : (-12'h14)) ? $unsigned(w100) : (-26'h16))) ? (^w80) : $unsigned((-24'h2)));
assign w38 = $signed((~|(((w46 == w74) < ((-20'h1e) ? w44 : w62)) ^ (29'h13))));
assign w39 = w91;
assign w40 = {($unsigned((10'h10)) >= ((-12'h4) ? w42 : w75)), ((w76 ? w69 : (-18'hf)) - $unsigned((-8'h2))), ($unsigned(w58) >= $unsigned(w99)), $unsigned({(6'h1b)}), $signed((|(19'h4))), $signed((w81 !== w56)), (|(-7'he)), w72, $signed(w70), (^~w81), ($signed(w61) < (w95 ? (-28'h0) : w62)), (^~(w1 === (-3'h1a))), (+{(-14'h1c), w66, w4, (-8'h19), w48, (25'hd), (9'h2), w45, w52, (-17'h14), (-18'h1b), (-18'h11), w93, (17'hc)}), $unsigned((10'hd)), ({w46, w7, (-11'h18), (21'hc), (-28'h6), (-23'h1a), (-18'h13), (-19'h6), w78, (-25'h1), (8'ha), w49, (-9'h19), w60, (-23'hc)} ? (w58 ? (-28'h14) : (22'h12)) : (w87 <= (13'h4))), ((w44 != (-2'h17)) ? (-21'h4) : ((-7'h7) ^ w3)), (~&$unsigned((11'h17))), w47, (^(4'h15)), $unsigned((w90 ? w77 : (16'hd))), $signed((w84 ? (1'h1a) : (-7'hc))), ((-w63) ^~ w45), (((29'h10) | (14'h15)) ? (24'h11) : (^w49)), ({(-4'h15), (6'h1b), w46, (-29'hd), (-9'h1), w2, w60, w53, (29'h2), (-20'h4), (-4'h11), w66, (20'h15), w8, w60, (-30'h18), w78, (32'h11), (-1'hc), w57, (15'hb), (-5'he), (-5'h16), w89, (28'h12), w6, w59, w1, (-25'he), (11'hf)} ? (w95 ? w77 : (19'h1)) : $unsigned(w44)), w62, (w54 - (~&(-13'h1d))), $signed((|(-1'h7))), ({w45, (35'h1d), (2'h8), (13'h13), (27'h1c), (-27'h11), w80, w78, (25'ha), w92, (19'h14), w63, w94, w47, (-14'h1e), (-1'h1b), w94, w49, w5, (-5'h4), (-16'hc), w90, w76, w49, (26'h19), (-13'h19), (-23'h19), w47, w52, (-9'h5)} === w66), (8'h11), $signed(w54)};
assign w41 = (w76 ? ((({w48, (-17'h0), (-10'h1c)} == (w53 != (23'h1b))) > (^~$unsigned(w93))) >= ((w74 || (31'h4)) ? (w64 ? w6 : (27'h8)) : (-16'h17))) : ({(-19'hf), w72, w79, (15'h12), w62, (-3'hd), w89, w70, w60, w77, w63, (-11'h1d), w63, w48, w74} ? {(-22'h16), (-14'h1e), w83, w8, (18'h19), (-23'h18), (26'h14), w97, w77, (23'h10), (23'h4), (-13'h1e), w95, w53, (3'h11), (-19'hc), (-3'h3), w44, (-5'hd), w69, (6'h14), (18'h6), (-30'hc), w96, (-15'h12), (-27'h1), (-19'hc), (-9'h12)} : {(13'h3), (24'h1a), (23'h1), (1'h4), w45, w50, (-34'h14), (24'h14), (-34'h1d), (7'h1c), (-18'h1d), w71, (-15'h7), (-16'hf), w45, (2'hd), w43, (13'h15), (11'h11), (-23'h0)}));
assign w42 = ((|{(29'hf), (-33'ha), w90, (14'h19), (7'h1b), (12'h18), (23'h12), w75, (-14'h17), w7, (20'h1a), (-19'hb)}) != (~&(-1'h15)));
assign w43 = (|($unsigned($signed((w1 ? (9'h7) : (-3'h19)))) << {(27'h2), w2, (-5'h16), w46, w2, w53, w7, w87, w68, w53}));
assign w44 = $signed(w67);
assign w45 = $unsigned((~^((~&(~&(-27'hc))) ? (w71 - {(27'h13), w72, w7, (24'h9), w61, w90, (-20'h7), w46, (-26'h15), w70, w87, (13'h1d), (14'h1a), w91, (-13'h5), w81, w1, w60, w62, (-27'hd), (6'h9), w57, (5'h18)}) : (-$unsigned((-22'h13))))));
assign w46 = ($signed(((11'h9) ^~ $unsigned({w90, w69, w75, w54, w96, w87, (26'h19), (-32'h1), (5'hf), w47, (1'h6), w6, w66, w6, (-27'hb)}))) ? w64 : {(w10 > w71), ((6'h1d) >= w77), {w1, (-27'h2), w70, (23'h10), (30'h10), (22'h13), (-22'h11), (-16'hb), w47, w10, w62, w52, (-28'h14), (-18'h12), w80, w53, (10'h15), (8'h5), w52, (21'h6), (26'h3), (26'h10), w76, w10, w72, w59, (-10'h2), w90, w73}, w99, ((-23'h15) ? (-30'h3) : (-15'h3)), (11'h5), (w64 ? (-9'hb) : w63), (-28'h1d), $unsigned(w59), ((15'h1b) || w7), {w49, w90, (-4'h18), w5, w10, (1'h5), w80, w80, (13'h3), w96, (-4'h18), w98, w99, w73, (-4'h1d), (8'h8), w97, (18'hc), w70, (18'h3), (23'h3)}});
assign w47 = (22'h9);
assign w48 = {w95, (^~(21'h12)), (-23'h1d), (((-13'h12) ? w6 : w89) ? (w86 ? (24'h18) : (-5'h9)) : (28'h5)), ((w97 ~^ (33'hd)) ? ((24'ha) < w87) : (6'h1c)), {(-10'he), (-29'hf), (32'h11), (-20'hf), (-26'h11), w99, (-8'h1b), (19'h6), (-19'h1e), (20'h18), (26'h18), w85}, (-19'h19), w90, w86};
assign w49 = (^{(8'h13), ((16'h8) < w85), (|(11'h1d)), ((31'h1e) ? w88 : (-30'h12)), (|(-22'h12)), (^w57), (w69 ? (21'h1c) : w58), (w96 << w64), $signed(w61), $signed((16'h19)), {(-8'h1), (-4'h8), w92, (-6'h7), (-22'h15), w78, (5'h16)}, (&(30'hc)), (w58 === w91), (~^(-11'h9)), (18'h5), w1, {(17'h1b), (-29'h18), (29'he), (-13'ha), (9'h1e), (-11'ha), (26'h2), w76, w96, w63, w73, w78, (-4'h0), (27'h18), w63, (14'h5), w77, w99, w82, w50, (-7'h1e), w80, (3'h10), w50, (7'h18)}, (8'h6), ((-4'h15) << w50), (w73 >= w65), (-29'h2), ((8'h9) ? w76 : w59), (-20'h11), {(-2'hf), w1, (11'ha), (19'h1b)}, (19'h19), $signed((8'h5)), (17'h1), $unsigned(w3), ((14'h1c) * w97)});
assign w50 = (($signed({w98, w86, w56, w64, (-24'h5), w51, (-8'ha), (-4'h10), (-27'h9), (29'h13)}) <<< $unsigned({w61, (17'h12), (16'h1d), (2'h8), w80, (-30'hb), w84, w8, (-8'h16), (-13'hd), w83, w67, w61, (-28'h1), (8'h10), w100, w98, w83, (-27'h18), w63, w88, w71, w81, (24'he), (-3'h8), w76, (25'h7), (18'h1a), w9, (-2'hc)})) ~^ {(-w97), (&(-26'hd)), (w2 === (13'hb)), (~^(26'hd))});
assign w51 = $unsigned($unsigned($unsigned((&$signed((-19'h13))))));
assign w52 = {{w63, (27'h18), w99, (-24'h9), w71, (-18'h7), (5'h15), w3, w89, w85, (17'h13), (14'h16), w64, w78, (-6'he), (1'h9), w97, (30'h1e), w75, w55, (-14'h1), (-13'h1c), w72, (-25'h15), w77, (-2'h1d), w54, w78}, (20'h1), (-13'h6), ($signed((-30'h10)) ? (w80 >> w70) : {(-29'hf), (12'hf), (-16'h1), (25'hd), (34'h18), (11'h9), w73, (-29'h1), w81, (-17'h1a), (-29'h5), (-6'h0), (-10'h8), (-25'h1d), (12'h11), w3, (15'hc), (-8'h18), (-1'h11), w86, (-25'h19), w10, (-13'h18), (17'hc), (-21'h19), w91, w89, (-30'h7), (-17'h14), w55}), $signed((2'hd)), $unsigned(w74), $unsigned($signed((1'h6))), w71, ((-10'h9) ? (|w87) : (26'h8)), (-$signed(w65)), w60, w94, (16'h16), w79, ((27'h15) ? (w98 ^ (20'h14)) : w55), $signed(((17'h17) ? w55 : w71)), (-22'h9)};
assign w53 = ($signed({(9'h2), w87, w6, w96, (22'hb), (-28'h1b), w69, (-23'h5), w59, w100, w95, (-26'h16), w95, (-12'h1c), (-20'hc)}) ? (-19'h1) : ((w95 ? $unsigned(w92) : w81) | $unsigned(((w78 & (-17'h1e)) !== {(-9'h17), w1, (15'h4), (-25'h3), w95, (-20'h1b), (9'hb), w81, w5, (29'h13), (-13'h8)}))));
assign w54 = $unsigned(((-28'h7) ? (((22'hf) > (-7'h11)) ? w93 : (~&(-21'h18))) : {w59, (-16'h10), (-1'h5), w86, w62, w4, (10'h3), (-17'h16), w56, w96, (-17'h14), (-28'h8), (27'h19), (-29'h12), w56}));
assign w55 = w85;
assign w56 = ({(^w72), (~&(-27'h8)), (+(-22'h3)), (&w94), w69, (w96 ^~ (23'ha)), (~|w76), $signed((-10'h2)), (~|w2), ((-4'h1d) ? (30'h16) : w67), (-29'h4), $signed(w57), (w94 && (-24'h1)), ((-22'h7) <= (6'h18)), w92, w71} * $signed((((-21'h12) ? (-21'h15) : w5) ? (^(w75 ? w70 : w6)) : (12'h1c))));
assign w57 = (-4'h14);
assign w58 = (3'hd);
assign w59 = $unsigned({(-11'hb), w8, (w76 ? w82 : (-29'h16)), w86, (w4 ^ w62), {(-22'h16), (-12'h9), w7, w81, (-17'h0), w81, (-1'h1e), w65, w67, w90, w10, w96, (-11'h19), (-7'hb), w93, (3'h8), w9}, ((26'h1b) ? (4'h1a) : (-30'ha)), ((-31'h10) >= (-18'h1b)), $signed(w82)});
assign w60 = w77;
assign w61 = ({w68, (^~w74), {w67, (19'h2), w3, (7'h9), (17'h5), (-22'h17), (13'hb), (-2'hb), w95, w72, (15'h2), w82, w65, (14'h12), (-18'he), (-10'h12), w71, w69, w82, (8'h11), w78, w98}, w96, $unsigned(w67), {w79, (13'h6), (22'h17), (-28'h17), w100, w70, (19'h1c), (12'h9), (15'h13), w82, (-14'h4), w85, (27'h9), (-8'h1c), w63, w10, (-19'h1d), w86, w93, (31'h7), (-23'h4), (34'h1), (5'h12), w63, w91, (10'hf), (30'h1c), w2, w64, (-5'h16)}, (w97 ? w81 : w3), {w91}, (w100 ? (-17'h6) : (7'h6)), ((-8'ha) ? (20'h2) : w7), {(-29'h4), w64}, (-(-10'h2)), {(-17'h1a), (-28'h1b), (-13'h5), (-26'h16), (-23'h1a), (-11'h1c), w10, (12'h1d), w10, (19'h17), (-22'h1a), w6, (15'ha), w4, w93, w81, w100, w100, (-16'h2), (12'h13), w75, w4, w77, (4'h1)}, {(-16'h8), w64, w74, w83, w87, w87, (24'h1d), (-18'h19), w83, w9, w97, (-12'h0), w75, w94, (-19'hb), w70, (1'h1a), w94, (30'h1b), (4'h2), (-32'hd), (5'h2), w2, w83, w68, w7, (31'h1a), w79, w65}, {(16'h5), (-1'h12), (-13'h4), w91, (-8'h0), (-18'h1e), w75, w74, w10, (3'h14), (-4'h19), w89, (-15'h7), (26'h8), w84}, ((-6'hc) ? (-5'h1b) : w5), $signed(w88), $signed((-3'ha)), (w84 + w90), {w87, w6, (-25'h1e), w5, (27'h3), w67, w70, (24'h11), (20'hc), (21'h15), w74}} ? w64 : {(w7 > w67)});
assign w62 = {{(-23'h4), w91, (-15'h4)}, w98, ((|w75) << ((-6'hd) == (12'h1c))), (23'hb), ((16'hc) | $unsigned(w3)), w77, (w5 ? $unsigned((-5'h1d)) : (18'hf)), ((-w82) ? ((4'h1d) || w1) : ((6'ha) ^ (20'hf))), w8, (-17'h11), ({(-21'he), w96, w67, w79, (3'h11), w73, w70, w94, w6, w89, (-27'h1), (25'h14), w68, w7, w91, (-21'h19), w63, w63, w99, (18'h7), (-26'h1), w100} - (11'h1b)), (((-26'h14) * w7) * (w8 !== (-23'h14))), {w8, (-6'h1a), w84, w69, w64, w75, w91, w71, w88, (21'h16), (-30'h15), (14'h15), (26'hd), w86, (16'hb), w8, w80, (29'hb), w93, (15'h10), (27'h12), (3'ha), w10}, (((5'h4) && (-29'he)) + w10), (w63 < (-12'h1)), $signed({w79, (26'h13), w75, w7, w79, w71, (8'h1), w88, (24'h2), w86, w63, (-30'h1c)}), {(-15'h14), w6, w97, (-17'h1c), (-6'h5), w98, (12'h3), (23'h17), w73, w66, (17'h12), (-8'h3), (9'h17), (-15'h15), (8'he), w9, (-13'h0), (18'h6), (-17'hb), w83, (4'h19), (19'h1a), w83, (-6'h5), (8'h18)}, (^((-22'h18) ? w63 : (24'h1a))), ($signed(w68) ? w2 : {w73, (-16'h13), w78, w78, w82, w65, w84, w90, w66, w1, (-28'h1e), w100, (-27'h5), w77, (-8'h1d), (-12'h13), w99, w3, w3, w95, (29'h18), (-19'h3), w81}), (19'h2), {w88, w91, (2'h8), w65, w93, (23'h11), w2, (-22'h18), w87, w91, (-27'ha), w77, w71, (5'h1e), w70, (-3'h12), (9'hc), w86, (-11'h3), (28'h19), w9, w77, w70, (-18'h15), w72, w74}};
assign w63 = {((|w65) ? (w8 * w77) : (8'h12)), (^(~^w8)), ((~&(21'h1e)) & $unsigned((-31'h6))), (13'h13), {(8'h8), w95, (14'h2), (10'h6), (25'h1a), w71, w94, w99, w88, w72}, (-3'h15), (w1 || (w94 ? (-5'h1) : (-13'h16))), ((-1'h8) * (^w72)), w78, $signed((~|w10)), (w94 !== $signed(w8)), w75, $unsigned((w6 ^~ (-10'h12))), (^~{w100, w10, (15'h16), (25'h8), (3'hd), w4, w96, (22'he), (9'h10), (3'h2), w99, (-12'h11)}), {w4, (-4'h1c), (11'h10), w74, w83}, w85, ((~|(-3'h7)) ? (16'h17) : {w86, w80, (18'h1), w75, w94, w7, (5'h7), (32'h15), w77, (-7'h9), (-30'h8), w88, (-6'h5), w66, w1, (-27'h9), w71, (29'h14), (14'h12), w98, w10, (20'he), (-16'h19), w83, w80, w74, w72, w9})};
assign w64 = (w94 ? (w82 ? w67 : (-7'h9)) : (^~$signed((+((14'h16) ? w81 : (-13'h15))))));
assign w65 = ($unsigned($unsigned({(13'h4), w79, (20'he), w91, (10'hb)})) ? {w72, ((19'h4) ? (25'h19) : (-22'h0)), ((-31'h6) ? (15'h9) : (21'h18)), ((-4'h17) ? (20'hb) : (6'h1e)), w7, {(-12'h18), (27'h1c), w86, (16'h18), w89, (-12'h0), w84, (-19'ha), (28'h13), (-19'h15), (-11'h17), (2'h1b), (-22'h7), w76, (15'h9), w88, (24'he), (16'h5), (-4'h1b), w71}, (-27'h1b), (^~w96), ((-12'h2) ? (24'h19) : w73), ((25'h2) ? w100 : w66), {w96, (-28'hd), w72, w98, w98, w3, (-7'h14), w66, w94, w80, (-17'hd), w95, (-26'he), (23'hc), w90, (-7'h18), (29'h11), w6, (30'h10), w72, w92, w3, w72}, ((-20'h1) ? w94 : w1), $signed(w77), {w2, w75, (9'h16)}, w84} : ((-22'h1d) << w84));
assign w66 = (^~w96);
assign w67 = (w6 + $unsigned((|({w76, w85, (-29'h5), (-18'h12), (4'h14), (23'h19), (1'h1e), w80, (18'hb), w1, (4'h3), w73, (-13'hc), (18'h1), w5, w100, (-6'h7), (-7'h13), w6, w74, w95, w79, w87, (28'h9), w83, (-4'h4)} >> $unsigned((-29'h1a))))));
assign w68 = (~&$signed(w3));
assign w69 = (~^(!($unsigned(w9) - w8)));
assign w70 = w2;
assign w71 = ((-26'h1a) ? $unsigned({(-15'h6), w98, w82, w86, w8, (8'h14), w88, w86, (11'h1b)}) : {(w8 ~^ w92)});
assign w72 = {(27'h14), w10, (((-28'h11) <= (9'h16)) ~^ $unsigned((-5'h6))), (21'h13), ({(15'h9), w8, w80, (-28'h5)} & $unsigned((-2'h13))), (-$unsigned(w75)), ((w87 ? (-15'h2) : (-7'h1e)) ? $unsigned(w75) : $signed((-11'h9))), (~^w88), (14'h15), (!(-13'he)), {(5'h10), w85}, (~|w94), {(20'h15), w94, (-20'hb), w93, (7'h7), (28'h13), (-26'h10), (-16'h7), w80, (-17'hf), (21'he), (2'h13), w90, w97, w74, w87, w6, (-14'he), w95, (-20'ha), w76, w73, w8, w88}, (~&$unsigned(w98))};
assign w73 = ((-4'hf) ? {(~&w3), $unsigned((-28'h17))} : (w8 << (8'h17)));
assign w74 = (32'h1c);
assign w75 = (~&w81);
assign w76 = {(w92 * $signed((-17'h6))), ((w5 ? (24'h5) : w86) ? (~|w6) : w95), ((w91 <= w93) + (w6 ? w88 : (-10'h4))), ($unsigned((15'h5)) << {w2, (-14'h1c), (-9'hf), (-22'h3), w82, (9'h1), (-11'h1), (25'h14), w91, w79, w87, w97, (-26'h18), (23'h2), w92, w3, w1}), w83, ($signed((21'h3)) === {(-10'h11), (-2'h1c), w5, (11'h4), (-22'h11), w93, (-16'h5), (-1'h9), w90, (-13'h1), w86, w87, (12'h3), (-22'h8), (28'h18), (-28'h18), (-20'h14), w100}), (((-22'h11) >= w93) ? (-23'hd) : (-(23'h1))), $unsigned(w5), ({(5'h6), w81, w90, w83, (-30'h1e), w98, w85, (-18'h11), (-6'h2), w4, (-7'h14), w77, w88, (8'h1b), w90, w100, w1} ? ((-18'he) ? (-19'h7) : w91) : {(-28'h18), w94, (-7'h1), (16'h4), w3, (-8'h10), w7, w8, w5, (-18'h5), w94, w78, w10, (23'ha)}), (w80 >>> (-5'h12)), (&w2), {w7, w79, w86, w84, (-7'h11), w2, (-1'h10), w2, (25'h2), w99, (-13'h1b), w3, w100, w87, w86, w91}, ((w88 ? (-19'h4) : (-14'h3)) - w99), (14'h17), {(-10'h7), w85, w95, (2'h11), (-16'h9), (12'h7), w6, (16'h19)}, ((6'h1b) ^ (&(22'h16))), {(-3'h1), (-10'h9), (-5'h12), (-18'he), (27'h19), w96, w88, (8'h11), (-23'h0), w85, w4}, (~&{(-26'h1), w80, w99, (22'h8), (1'h10), (-24'h15), (-27'h1a), w88, (-19'he), w5, w80, w92, w85, (19'h9), (21'h4), w89, (-13'h10), (-28'h7), (-6'hf), (8'h19), (23'h11), (-3'h3), w87, w78, (17'h1d), w99, (4'h14)})};
assign w77 = {$unsigned((~^w88)), (13'ha), ((w3 <<< w98) ? $unsigned(w96) : w1), (-10'h1e), $unsigned({w96, (-28'h8), (4'h1c), w8, (16'h1), (-9'h5), w97, w5, (-15'h1d), w99, (-15'h3), (17'h14), (-29'he), w4, (-26'h1), (18'ha), (31'h10), (-4'hf), (-29'hf), w86, w92, w89, w91}), (&{w83, (-5'hb), w95, w2, (-32'h19), (-15'h3), (-12'hd), w93, (4'h13)}), {(14'h18)}, (-27'h18), {w84, (-25'h13), (30'h18), w79, (-15'h13), (13'h16), (-23'hc), (-5'hc), (9'h5), (20'h14), w89, w100, w97, w4, w3, (-23'h16), w9, (-33'h3), (3'h3), (-12'h7), (18'h14), (-2'he), (-2'h0), w78, w80, w7, w99, w88, (-11'h19), (-30'h19)}, {(-23'h16), w91, (-1'h1b), (-24'hb), (-18'h10), (-32'h5), (24'h6), w87, (-10'h17), (23'h19), (-1'h3), (16'h13), w98, w83}, {w86, (12'h1c), w95, (14'h8), (-5'h19), (17'h1e)}, {w84, (-7'h3), (-20'h13), w91, w83, (20'h10), w78, (-26'h17), w81, (-1'h11), (-28'h19), (-9'h8), w100, w84, w83, (-12'h17), w85, w6, w100, (-4'he), (25'hd), (-16'he), (16'h18), (-25'h10), (-3'h18), w97}, ((w8 ? w8 : (-8'h9)) || $signed((-19'h4))), {(-1'he), (-23'h9), (-24'hd), w85, w4, w10, (18'h1a), w91, w3}, ((29'h1c) ~^ w86), {(-11'hc), (-7'ha), (26'h5), w83, (-23'h1e), (-25'h7), w82, w98, w98, w90, (-7'h7), w87, w94, w95, w1, w87, w79, w87, w81, (-23'h17), (13'h8), (-10'h0), (-30'h8), (26'ha), (-14'h1a), w98, w81, (23'hc)}, (~&((-30'h1c) ? w6 : w6)), ({w87, (22'hb)} ^~ (w5 ? w85 : (-17'h18))), (w79 !== w100), $unsigned(((1'ha) < (4'h16))), (((-12'h3) ? (-10'h19) : (21'h1c)) == ((30'h1d) ? (-17'he) : w6)), (((-19'h1b) ? w85 : w87) ^ (-29'h11)), ({w88, w90, w5, w2, w89, (-18'h1b), w92, (-27'h1), w6, (25'h1), w1, w85, w1, (-8'h15), (-28'hc), (-8'h0), w87, w92, w95, (-4'h6), (-30'hb)} ? {w81, w78, (11'h2), w8, w1, (1'h15), w8, w5, (5'h7), w100, w86, (-2'h10), w5, (-32'h7), w96, w98, w91, w2, w100, (21'h1e), (-29'h6), (16'hd), w3, w83} : (|w6)), {(-1'h14), (-17'h13), w80, w10, (-5'h7), (4'h16), w83}, {(21'h6), w99, (30'h13), w96, (6'h10), w88, w99, (-18'h12), (7'h11), (-6'h1d), w94, w80, w99, (-22'h11), w99, w84, w94, (16'h7), (7'h4), (-3'h5)}, (-(w87 ? w10 : w88)), ({w83, w6, w94, (-19'h19), (-21'h15), (-19'h0), w97, (-27'h19), (9'h5), (-4'h0), (22'h13), w99, (6'h11), (-26'hd), (23'h11), w9, (-6'h7), (-16'h1a), (22'h1b), (-12'h8), w89, (7'h1d), (33'h19), w94, (29'h1b), w1, (-2'h18), (10'he), (29'h19), (-28'h7)} ? ((-28'h1a) * (4'h8)) : {w85, w91, (-20'h12), (4'h1c), (-19'h3)})};
assign w78 = (~&(^((18'h1) - ((-12'h2) ~^ {(-8'h1b), w82, (29'h13), w88, w5, (14'ha), w96, w93, (-21'h0), w3, (28'h3), w5, (23'hc), (-19'h7), w9, w10, (16'hb), (-8'h11), (25'h8), (15'h3), (3'h2)}))));
assign w79 = ($signed((|{(-13'h1c), w93, (-10'h1b), (-24'h13), (4'h1c), (30'h1d), (4'h19), (-18'h6), w6, w92, w10, w4, (11'h2), (-7'h6), w90, w5})) ? (-15'h2) : (~^((-13'h18) <= ((-1'h1d) >= (w80 ? w2 : (-20'h1))))));
assign w80 = ((-18'h3) ? ($signed((&(-2'he))) ? ((-14'hc) ? (^~(30'hc)) : (~|(-24'ha))) : ({(21'hf), w93, w7, w83, w88, (-4'h16), w89, (-25'h15), w96, w94} || w85)) : $unsigned($unsigned(($signed(w3) * (-w9)))));
assign w81 = (-9'he);
assign w82 = {$unsigned(w7), ((&w97) ? $signed(w86) : (w6 > w99)), $unsigned((-w6)), (+w84), w3, ((+(-14'h14)) ? ((-5'hf) ? w1 : w95) : ((-4'h14) === w92)), (!((-27'ha) ? (-10'h2) : (16'h4))), (((28'h1e) | w87) ? (w86 === (33'hd)) : ((3'h1c) & w7)), (((-19'h4) ? (-11'h14) : (15'hd)) ? {w9, (-25'hb), w90, w93, (-10'h7), (-5'h12), w86, w98, w95, (27'h1b), (-18'hc), w87, w5, (4'hf), w84, w6, (30'h1c), (27'h11), w88, w89, w88, (-3'h10), w4, (12'h19), (-21'hb)} : w83), (^~$unsigned((-8'h12))), {w96, w92, (25'h5), (-24'h6), w85, w87, (24'h2), (-27'h1d), w84, (28'h1b), w95, w9, w84, (27'h6), (-7'h1e), (-25'h8), w91, w3, w89, w97, (-16'h16), (-5'h8), (-30'h14), (-23'h10), w5, w88}};
assign w83 = $unsigned({(-15'h1e), w96, (~&(6'hc)), {w84, (29'h17), w84, w97, w88, (-26'h1e), (29'h1e), (9'h19), (28'h1b), (25'h1b), (-5'h1b), w96, w86, (11'h1b), (22'h12), (26'h5), w93}, (16'h16), (-w1), {(6'h13), (28'h5)}, w2, w4, {w95, (-25'h1e), w3, (5'h9), w92, w94, w86, (4'h2), (11'h14), w7, w7, w3, (19'ha), (-26'he), w88, (17'h1e), (-11'h14), w2, w99, w6, (-23'h15), w85, (13'h14), w89, (4'hb), w4, (-16'ha), w90}, $signed(w94), (w98 >= (-13'hc)), (w91 ? w6 : w93), {w10, w9, (3'h11), w8, w92, (3'h10), (-12'h1c), w93, w94, (10'h1e), w4, (3'h18), (-2'h14), (-26'h6), w92, w8, (-4'h14), w84, w94, w90, (30'h7)}, ((-3'h8) ? (-12'h15) : (-6'h18)), (w100 ? (8'h3) : (23'h6)), $unsigned(w88), w8, ((3'h10) ? (23'h5) : (-17'he)), (20'h5), $signed((-26'h4)), {w94, w7, w99, (7'h10)}, {w85, w1, (-15'h1b), (8'h12), (-16'h7), w10, (17'h14), (-24'h10), w84, w88, w99, (-25'h19), (-20'h9), w98, w84, w99, (-16'h1b), w90, (3'h16), w7, (22'h16), (12'h3), w100, w100, (-5'h1a), (-6'h6), w3}, ((19'h1d) ? w6 : (32'h8)), (30'h1c), ((22'h1d) ^~ (26'h1c))});
assign w84 = w92;
assign w85 = w10;
assign w86 = (8'hc);
assign w87 = (^~$signed((({w100, w90, (23'h5), w6, (-4'h16), w92} ~^ {w88, w93, (2'h10), w90, (-3'h15), w3, w2, w95}) ? ((4'hc) === $unsigned(w6)) : w100)));
assign w88 = {((-19'h1d) ? $unsigned((-16'h5)) : (-23'h9)), $unsigned({(14'h3), (4'hd), (-14'h1d), w95}), (!(-30'h14)), (-21'hb), (+(w1 ? w92 : w9)), (&(w96 - w5)), $signed(w2), ({w95, (-13'h1), (-29'h1d), (-18'ha), (12'he), w96, (2'h1c), (4'h15), w7, w10, w98, (5'h11), w4, w8, w95, (1'h6), w91, w6, w90, w96, w98, (23'h1)} && (w98 | w91)), {(7'he), w3, (9'h19), (-1'h8), (25'h18), w100, w4, (-20'h6)}, (~^(w10 ? (-7'h1c) : (-24'h15))), (-24'h18), $signed(w1), $signed(w91), (~&w10), ((-27'he) ? $unsigned(w89) : (13'h8)), w90, ((-20'h10) - (~&(-14'hd))), ((w92 >= w3) ? $unsigned(w94) : (^~(-12'h17))), $unsigned((w98 ? (-19'h5) : (11'h1c))), w92, w1, {w93, w2, (-29'h6), w89, (24'hf), w91}, (-18'hf), (-20'h12), {(30'hf), w1, w98, (-17'h0), w9, w98, (-14'h14), w5, w7, w100, w10}, $unsigned((^(4'h9)))};
assign w89 = (~^$signed($signed((7'h9))));
assign w90 = (w96 < {$signed(w1), {w4, w7, w8, (13'h10), (-13'hb), w95, w5, w91, (-6'h13), (-25'h1a), (30'h16)}, (w94 ? w98 : (14'h11)), (-(23'h1e)), w7, (^~(1'h16)), (w92 ? (1'h1b) : (8'h1d)), w96, (w1 ? (-20'he) : (-17'h16)), ((15'h3) ? (-24'h9) : (-8'h17)), w1, ((8'hf) != (-2'h1b)), ((-30'ha) ? (-21'h1) : (-2'h13)), w92, (!w8), (~^(-25'h9)), w6, (-7'ha), {w4, (-5'ha), w9, w96, w98, (4'h1a), w3, w8, w92, w98, w99, w99, (-2'h11), (20'he), w7, w10, w5, w97, w99, (-21'h1d), (-31'h6), w5, w5, (-10'h5), (-10'h8)}, (14'h13), {(-17'h7), w1, w93, (4'h8), w4, w8, (-15'h12), w94, (5'h1b), (-6'he), (14'hc), (-18'h13), w7, w97, (6'hb), (-24'h1b), w92, (6'h14), w6, (19'h5), (-5'h1e), (-28'h1), (28'hb), w98}, (~|(-16'hf)), ((-30'h2) & (19'hf)), $unsigned((21'h1d)), ((15'h6) ? (7'h4) : (30'h13)), $unsigned(w8), $unsigned(w6)});
assign w91 = (^~{(-10'h4), w92, (-11'h5), {w4, w1, (30'h10), (-13'h11), (-17'h17), w98, w93, w4, (16'h7), w2, (-9'h6), (21'h1c), (-21'h3), w1, (31'h1b), (19'h5), (-12'ha), w7, (22'h13), (-27'h19), (10'ha), (-1'hc), (-25'h1d), (25'h12), w7}, (~^(3'h11)), ((24'h4) ? w8 : (18'h9)), (|(-24'h19)), ((-7'hb) ? w2 : w92), (25'h3), w100, w4, ((-9'h10) ? w9 : (-3'h1c)), {(-9'hb), w6, (8'h17), (-10'h1d), w96, (-11'h15), (31'h7), (-20'h1a), w100, (-20'h1d), w92}, (~^w100), (+(-15'h18)), (w98 << (28'h7)), (~|(-10'h1d)), (23'h3), (w4 ? (17'h15) : w2), w96, w1, w96, w98, (w99 ? (-8'h9) : (-13'h1b)), w2, (9'h16), (~&(14'h5)), ((3'h9) < w3), ((1'hd) !== w6)});
assign w92 = (~&(~|w98));
assign w93 = $unsigned($signed(((w4 < ((-21'h8) & (14'h14))) ? (23'hf) : $unsigned(w5))));
assign w94 = ({{(32'h6), w1}, (~&w99), (w3 == (-15'h8)), ((-28'h17) ^ (6'h1)), (-6'h1), (w6 ? w4 : (-21'h10)), ((-9'h16) ? (25'h1d) : (-17'hd)), ((18'h1) > w97), (w4 > (6'h13)), (3'h8), (-17'h13), w96, w97, (^(-3'h4)), (^~w3), (6'h1a), {w1, w2, (-22'h19), w3, w9, w8, (12'h1), (26'h3), (8'h16), w8, (-21'h15), (9'h7), w95, w8, w100, (-15'h1e), (30'h14), w98, w10, w95, (-5'h3), w100, (12'h7), w95, w7, w4, (1'h5), (10'h3), w8, (27'h4)}, (w99 ? w96 : w100), (20'h10), (-12'h1c), w2, $signed((-9'h6)), (^~(32'h10)), ((-15'h8) & (-4'h5)), ((2'h6) ? w4 : w1), (-13'h4), w96} ? (&(-14'h1c)) : ((2'hb) | (~&(w2 ? w6 : (17'h16)))));
assign w95 = $unsigned(({w99, (-4'hf), w96, w7, (-6'h1), w8, (-2'he), (-7'h3), (20'h7), (16'h13), w98, w100, w100, w8, (26'ha), (23'h9), w7, w97, (-13'h17), w4, w5, w7, (8'h3), (33'h19)} ? $signed((~|w6)) : w96));
assign w96 = $signed({(|(-2'h5)), (^~w97), w98, (~&w3), (|w8), w4, (7'h14), {w5, (-13'h12), (4'h1d), w5, w6, (-31'h1a), w98, (30'h7), (-18'h1c), w5, w3, (-16'h1a), w1, w100, w3, w6, w3, (-30'h2), w8, (22'h1e), w98, (-24'h18), w4, w4, w7, w100, w10}, $signed(w9), {w8, w3, (10'h14), (31'h1e), w10, w100, (30'h12), (9'h7), w7, w10, (-6'h17), (-8'h0), (18'h4), (-18'h17), (-5'h1e), (6'h1), w9, w10, (28'h11), (18'h12), (-27'hb)}, ((-15'ha) ? w9 : w99), (w6 << w7), $signed((-23'h17)), (w2 * w3), (-w5), ((-1'h12) ^~ w97), (-(20'h1e))});
assign w97 = {$signed($signed((23'hd))), w2, {w3, w10, (-18'h3), (-9'h18), w8, w9, (-26'h5), (-19'hb), (25'hb), w3, (-24'h7), w6, (31'h6), (16'h14), (-6'h7), w10, w10, w8, (-30'h0), (8'h10), (-6'h8), w7, (-18'h15), w98, (-15'h11)}, $unsigned((w9 ^~ (21'h1d))), ((^(-22'h15)) ^~ w2), (^(w10 ? w2 : w98)), (w5 ^ $unsigned(w6)), {w6, (28'hd), w100, w2, w98, w7, (2'h17), w9, (-32'hf), (-20'h19), w4}, ((w7 !== (-18'hf)) >> $signed(w6)), $signed((+w9)), {(36'h8), w99, w5, w10}, ((-18'h13) ? (w100 ? (-15'he) : (-20'h6)) : (~^(-24'h9))), {(-24'h11)}, ((-(-5'h14)) <= (~|(19'h19))), (19'h5), (-14'h10), ($signed((18'h6)) >>> ((13'h14) ? w6 : (-16'h10))), $unsigned(((18'h1e) != w8)), w10, (w1 === $signed(w4)), {w10, w1, w10, (-19'he), (-21'h0), (-5'h13), (3'h1c), w100, (24'hc), (-4'h0), (-28'h6)}, ({(24'hb), w7, (27'h7), (16'h19), w4, (-11'h13), (2'h1d), (-13'h10), (6'h10), w98, (-18'h16), w98, (-30'h5), (17'h10), w6, (-23'h11), w3, (-15'h6), (29'h1b), w3, w10, (3'h6), (3'h7), (15'h1b), w3, (-12'h6), w2, (-25'h1e)} ? $unsigned(w10) : {w3, w1}), {w8, w5, w2, w9, (-10'ha), w99, w98, (28'h1), w3, w3, w2, w6, (14'h3)}, (w4 ? (!w8) : ((-7'h1c) * w5))};
assign w98 = (3'h3);
assign w99 = (({(2'ha), w100, w3, (7'he), (22'h10), w5, w6, (16'h9), w9, w1, w1} !== $signed(({w6, w6, (-18'ha), w1, w7, (-1'h3), w6, w5, (16'h19), w100, (-4'h16)} && ((-16'h18) ? (16'h18) : (30'h1a))))) ? {(&(-18'h13)), (25'hb)} : ($signed($unsigned((7'ha))) ? w2 : (15'h18)));
assign w100 = (~^(22'h11));
assign y = {w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100};
endmodule
