module test_module(y, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10);
output wire [1393:0] y;
input wire [8:0] w1;
input wire [25:0] w2;
input wire [24:0] w3;
input wire [16:0] w4;
input wire [29:0] w5;
input wire [28:0] w6;
input wire [21:0] w7;
input wire [22:0] w8;
input wire [29:0] w9;
input wire [20:0] w10;
wire [18:0] w11;
wire [2:0] w12;
wire [18:0] w13;
wire [17:0] w14;
wire [28:0] w15;
wire [28:0] w16;
wire [12:0] w17;
wire [21:0] w18;
wire [8:0] w19;
wire [20:0] w20;
wire [16:0] w21;
wire [10:0] w22;
wire [15:0] w23;
wire [26:0] w24;
wire w25;
wire [1:0] w26;
wire [1:0] w27;
wire [25:0] w28;
wire [24:0] w29;
wire [1:0] w30;
wire [13:0] w31;
wire [18:0] w32;
wire [25:0] w33;
wire [23:0] w34;
wire [24:0] w35;
wire [25:0] w36;
wire [26:0] w37;
wire [4:0] w38;
wire [26:0] w39;
wire [21:0] w40;
wire [2:0] w41;
wire [6:0] w42;
wire [21:0] w43;
wire [12:0] w44;
wire [1:0] w45;
wire [2:0] w46;
wire [2:0] w47;
wire [13:0] w48;
wire [10:0] w49;
wire [25:0] w50;
wire [19:0] w51;
wire [4:0] w52;
wire [11:0] w53;
wire [17:0] w54;
wire [20:0] w55;
wire [18:0] w56;
wire [22:0] w57;
wire [22:0] w58;
wire [15:0] w59;
wire [3:0] w60;
wire [24:0] w61;
wire [9:0] w62;
wire [6:0] w63;
wire [17:0] w64;
wire [22:0] w65;
wire [8:0] w66;
wire [23:0] w67;
wire [17:0] w68;
wire [6:0] w69;
wire [9:0] w70;
wire [23:0] w71;
wire [13:0] w72;
wire [16:0] w73;
wire [11:0] w74;
wire [24:0] w75;
wire [24:0] w76;
wire [15:0] w77;
wire [13:0] w78;
wire [16:0] w79;
wire [4:0] w80;
wire [5:0] w81;
wire [14:0] w82;
wire w83;
wire [28:0] w84;
wire [7:0] w85;
wire w86;
wire [17:0] w87;
wire [1:0] w88;
wire [22:0] w89;
wire [2:0] w90;
wire [25:0] w91;
wire [25:0] w92;
wire [7:0] w93;
wire [25:0] w94;
wire [7:0] w95;
wire [5:0] w96;
wire [29:0] w97;
wire [7:0] w98;
wire [24:0] w99;
wire [14:0] w100;
assign w11 = $signed((-29'h9));
assign w12 = $signed($signed((-18'h7)));
assign w13 = {((w60 | (27'h9)) ? {(27'h1c), (-27'h1c), (-7'h18), (13'h15), w59, w48, w54, (8'h4), w18, (-2'h1c), (-17'h5), w78, w31} : (-8'hc)), {w97, w60, w23, w87, (-20'h7), (-19'hb), (-9'h2), (-15'h4), w33, w30, w49, w27, (29'h2), w41, (-8'h18), w55, w26, (19'he), (-10'h15), w44, (14'h15), (22'h19), w24}, {(-22'h10), (-6'h14), w28, w75, w90, (-14'hd), w21, w92, w68}, w92, (-7'h1c), $signed((w23 || w14)), w3, w61, $signed((-4'h7)), w85, (-10'h3), ((^w54) !== $signed(w74)), $unsigned(((2'h9) ? w65 : (-19'h6))), w1, (~|(!w58)), (5'h15), (^(-19'h4)), ((w97 ? w61 : w61) && (w53 !== w3)), (+$signed((20'h1b))), w82, (((10'hd) ? (-3'h1a) : w4) > (+w16)), (11'hd), {(-13'h7), (28'hd), w62, w8, w42}, (w6 ? {(22'h9), w74, (-15'h1d), w18, w1, (22'h7), (-24'h8), w100} : {w60, (-28'h19), (17'h14), w67}), ((w16 >>> (30'h2)) ? (-30'h5) : ((30'h10) <<< (-11'hc))), ((~&(5'hf)) >> ((-6'h17) || w76))};
assign w14 = w30;
assign w15 = w46;
assign w16 = w42;
assign w17 = (23'h1);
assign w18 = ({$unsigned((-8'h1))} ? ({w73, (18'h2), (-17'h14), (-22'h1d), w6, w58, w48, w41, w43, (-2'hf), w100, (1'h9), w38, w74, w81, w89, w92, w23, w77, w37, (13'h6), (-23'h11), w60, w78, (-25'h1b)} ? (&((-7'h1d) ^~ w70)) : ({(15'h1), (22'ha), (-16'h3), (11'h10), (1'h1b), (-20'h10), (-13'h1b), (-23'h14), w48, (-4'h1a), w51, (-24'h1e), (-16'h18), w38, w30, w29, (-12'h5), w42, w44, w54, w20, (-4'h10), (27'h7), (3'h9), w73} ? ((-22'h18) ? (9'h1a) : (4'h13)) : (&(23'h1a)))) : (w79 ? $unsigned(((-29'h12) <<< (14'h4))) : (24'h10)));
assign w19 = ({(w71 | (22'h11)), w42, {(-23'h7), w7, w54, w26, w73, w54, (14'h1c), w32, w71, w52, w89, w2, w74, (24'h5), w6, w90, (19'h3), w91, (3'h8), w61, (-6'h1e), (31'hf), (-30'h11), (22'h1a), (-27'ha), (-35'he), w68, (14'he)}, {w86, (-25'h4), w51, w52, w38, (-3'h1), w60, (-3'h9), (28'h19), (-18'h13), (-22'h0), w20, (20'h15), w21, (-1'h5), w37, (29'h1e), w36, (-16'h10), (-5'h1e)}, $signed(w92), {w44, w29, w95, (-12'h3), w34, (-21'h2), w37, (-19'h7), (-21'h11), (-11'h10), (-11'h16), (-27'h13), (14'h1e), w34, (-22'h7), w59, (-12'h8), w57, (3'ha), w51, (23'h13), w89, w73, (24'h15), (-22'he), (17'h8)}, (|(-19'h8)), (w82 >= w51), (w39 ? (15'h1c) : w59)} << w91);
assign w20 = (~&{w31, (-1'h2), $signed((-11'h1e)), (~|(-10'h1d)), (w25 ? w80 : w44), $signed((-13'ha)), (-24'h16), (w55 ? w41 : w78), {w8, (21'h1a), w69, w34, w50, (14'hd), (5'hb), (-5'h11), (-2'h3), w28, w87, (-7'h1a), (1'hf), w83, (-22'h18), w72, w87, (-22'h14), (10'h1), (30'h10), w91, (-21'h19), w97}});
assign w21 = {(20'h6), {(-26'h1d), (-22'hc), w26, w33, w82, (-29'hb), w27, w72, (15'h12), w34, (-29'h8), w87, w40, (9'h9)}, ((w60 ^~ w65) ? (w99 ? (29'h17) : w41) : (30'h17)), ((w86 || w39) << (w22 ? w100 : (-4'h0))), {(13'he), w70, (-10'h13), w34, (20'h9), (24'hc), w76, w94, (13'h19), w95, w86, (-28'h16), (-9'h19), w87, (-29'h16), w96, w7, (-31'hd), (-24'hd), (18'h1d), w2, (27'hb), w80, (-4'hb), (27'h14), (8'h1c), w92, (-13'h14), (20'h8)}, ((-17'h1d) ~^ (^(12'h7))), $unsigned($unsigned((-23'h4))), {(-1'hb), (18'h5), (-25'h10), (-23'h5), w49, (28'hd), (25'h3), (18'h1d), w68, (27'h10), w9, (-15'h1), (17'h10), (24'h1c), (-4'he), w3, w2, w6, (18'hf), (-17'h1d)}, ($unsigned(w70) - (~|w58)), (^~{w43, (-16'h1d), w48, w48, w99, w68, w48, w99, w67, w93, w10}), {w28, (-22'h8), w80, w57, w37, w57, w73, (-30'h13), w45, (3'h1b), (9'h6), (-11'h8), (26'h7), (-6'h13), (16'h15), w56, (-25'h8), w81, (-4'h1a), (-20'h14), (28'h13), (20'h15)}, ((~|(15'h4)) ? {(19'h2), (-14'h1a), w46, w65, w42, w45, w4, w23, w36, (17'h14), (-28'ha), (-29'ha), (-5'h9), (-2'h8), w34, w30, (-15'h1a), w3, w2, w7, w29, w26, (-16'he), (22'h5), (-25'h7)} : (+w42)), ((~&(-3'h7)) | ((-15'h0) ? (-21'hd) : w34)), {w72, (-10'h1c), w28, w98, (-21'h19), w58, (-16'h12), (33'hf), (-12'h7), w96, (4'h2), w68, (3'h8), (25'h4), w65, (-11'h1e), (17'h5), w67, (26'h6), (31'h19), w47, w73}, (-(6'h11)), {(-8'h9), w72, w7, (-10'h1), w78}, (((8'h7) ? w9 : w72) ? {(-23'h18), w71, (-14'h3), w59, (2'hd), (-2'h3), w34, (-9'h1b), (26'hc), (-3'h1), (-24'h2), w55, (20'h4), w37, w7, w55, w77, w52, (-13'hd), w82, w10, w60, w63, (-12'h1)} : (12'h17)), w38, $signed($signed((22'h18))), {(-21'h1), (6'hd), w73, (23'h11), w47, w90}, w45, $signed({(-20'hc), w79, w87}), (~^(w54 || w6)), (w96 > (^(28'h16))), (~&{(6'hc), (-23'h1b)}), ($unsigned((30'h2)) ? (w53 ? w70 : (6'h19)) : (w57 ? w68 : (-7'h10))), (11'h15)};
assign w22 = ((12'h5) || (~^(16'h8)));
assign w23 = {{w40, w32, (-1'h16), (18'h18), (-19'h17), (-23'he), w41, w99, w33, w60, (-26'h1a), w70, (-10'h13)}, {w92, w87, (-7'h7), w59, (28'h1a), w98, w89, (27'h17), (-10'h5), (-16'h6), (11'hc), w52, w82, (7'hc), (6'h16)}, ($signed((-2'he)) & ((30'h5) + w8)), ({(12'h18), (22'hc), (13'h1d), (-24'h1c), w9, w1, (-6'h13), (19'h18), (-11'hd), w44, w42, (12'h1a), w33, w31, (-16'h3), (13'h15), w6, w67, (16'h3), w93, w10, (-2'h8), (15'hc), (16'h13), (-2'h8), (-25'h1d), (30'h3), w84, w55, (3'hf)} ? $signed((-31'h3)) : {w97, (-6'h6), w75, w52, w65, w98, (23'hb), w2, (-30'h1a), w4, (5'h16), (11'h2), w96, w67, (18'h3), w45, w10, w4, w58, w54, w100, w6, w83, (29'h1e), w49, w58, w68}), (-2'h10), (^(w1 >= (-27'h4))), (24'he), ((w58 << w42) ? (w35 - (-8'ha)) : (~&w7))};
assign w24 = ($signed((w94 << (-13'hc))) ^~ {(w57 ? (-19'h19) : (-22'h1b)), (w47 & (8'h12)), (w72 + w43), $unsigned((21'h18)), w4, $signed(w64), (+w26), (w45 ? (13'hf) : (-22'h10)), {w99, w2, w84, w38, w96, w99, w64, w52}, w32, ((29'h10) ? (-22'hb) : (30'h18))});
assign w25 = $unsigned($signed($signed((-5'h14))));
assign w26 = (12'ha);
assign w27 = (-3'h1c);
assign w28 = (-4'h5);
assign w29 = ((((19'ha) && ((18'h1a) ? w56 : w85)) ? (~&($unsigned(w99) ^~ {w39, (16'h10), w95, w43, (-20'h18), (-13'h3), w36, w48, (-21'hc), (-29'hf), w33, w87, w76, w84, w46, w83, (-1'h1e), (-22'hb), (-27'h13), (-12'hd), w49, w32})) : (6'h1e)) === $unsigned((32'h9)));
assign w30 = w7;
assign w31 = (26'hb);
assign w32 = (-11'h1c);
assign w33 = $signed({$unsigned((5'hb)), (w49 ^~ (18'h8)), w80, (-(21'h4)), (-(-19'h0)), (w90 ? w99 : (22'ha)), (w49 - (21'h7)), ((-2'h1) ? w46 : w69), (-15'h1), (w43 <= (2'h13)), ((-1'h15) >= (-21'h3)), (~|w1), (-3'he), $unsigned((-25'hb)), $signed((-4'h12)), $signed(w92), {w51, w72, w68, w87, (8'h18), (26'h8), (10'h12), (-10'hb), w82, w96, w52, w89, w99, w2, w62}, (w79 ^~ (-1'h11)), ((23'h1d) ? (4'h6) : w74), ((9'h1d) ? (6'hd) : (-1'h1d)), (w63 ? (29'h10) : (10'h6)), (w46 !== w99), (-24'h13), (w39 ? w93 : w60), (~^(20'h10)), {w73, w54, (13'hc), w35, w63, (8'hd), w52, w67, w36, w44, (4'h10), w77, w70, w64, w98, (-20'h1c), w4, w42, (22'hc), w52, w80, (14'h1), (-27'h1b), (-24'ha), w71, (16'h16)}, (w50 << (-26'he))});
assign w34 = {(-w2), ($signed((-15'h1c)) ? (w61 <= (31'h1e)) : (|w10)), {(6'h14), w79, w5, w1, w60, (13'h4), w38, (-28'hc), (-18'h16), w67, (6'h15), (-15'h1e), (25'h17), w41, (23'h2), (10'h19), (26'h15), (2'h6), w66, (-13'h1e), w87, w48, (16'h2), (26'hb), w53, w36, w98, (18'h1a), (-27'h9)}, (1'h1e), (((21'h19) !== w35) ? {(-4'h6), (-8'h12), w53, (13'h3), (-4'h1b), (-10'hb), w62, (26'h4), w99, (17'h2), (19'h8), (6'h7), w55, w93, (-21'h1c), w79, (-4'h5), (2'h1), (-3'h5), (-3'hd), w71, w61} : $signed(w46)), $unsigned(w60), w93, {(-17'h1a), (29'h1b), w73, w54, w66, w76, (15'h6), (-6'h15), (-18'h1a), w9, (-3'h1e), w38, (31'h7), w54, w46, w75}, ((~^w9) << w49), (-16'h1d), (~|{(-1'h19), (-21'h11), w92, (14'h2), (22'h18), w85, (5'h1c)}), $signed($unsigned(w86)), $signed($signed((18'h8))), (w77 ? (-10'h9) : w61), {w36, w40, w75, w83, (-29'h12), w90, w78, (18'hf), w48, (-26'h13), w69, w48, w41, (-37'hd), (-28'h1c), (6'h14), (-10'h1), (-16'h2), (-14'h7), (24'h14), (25'h10)}, w88, (-5'h1d), w58, $unsigned((-28'h2)), ({w41, (23'h1), (-12'h3), w92, w74, w57, (-14'h11), (34'h15), (17'h1a), w95, (24'h1e), (3'h17), w94, w67, w50, (-15'h18), (-11'h9), (4'h9), w89, (-8'h6), w6, w74, (14'he), w56, w56, (-16'h15)} <<< w6), ($signed(w81) | $unsigned(w5))};
assign w35 = $unsigned((~&$unsigned(({(-10'he), (1'h8), w91, (15'h1c), w74, (29'h1b), w68, w84, w79, w73, (30'h4), w53, (-11'h14), w83, (-19'h1d), (29'h4), w59, (-18'h10), w78} ? ((5'h1c) + (10'h5)) : (w62 ? (17'hc) : w36)))));
assign w36 = (((((-30'h1) || w51) ? w56 : (w85 > w40)) ? w70 : (w94 * w60)) * (32'h18));
assign w37 = $unsigned((-25'hd));
assign w38 = (((($signed((10'h11)) !== ((-11'h10) ? w50 : w82)) || $signed(w10)) | ((~&(-29'h1c)) ? ((-8'ha) ~^ (4'h15)) : $signed((-9'ha)))) ? {(w40 || w73), ((6'h6) ? (12'h10) : (-26'h1)), ((28'h1d) ? (25'hb) : (11'hd)), (|(25'hf)), w3, w51, (-31'h9), (w75 | w86), (-2'hd), (-25'h1e), (26'h1d), w40, (w95 <<< w51), (^w47), (-(19'h11))} : w40);
assign w39 = (~^({(23'h1c), w83, w45, w94, w94} ? (-31'hf) : ((-15'h8) ? $unsigned((18'h14)) : (w47 ? (39'h1c) : (-15'h17)))));
assign w40 = ({$signed((19'h12)), (-10'h9), $unsigned(w65), $unsigned((5'h15)), w73, w73, (24'hf), (w6 ? (9'hd) : (-5'hd)), $signed((10'h15)), w51, $unsigned(w4), (w5 + w60), (w4 <= w51), (w71 ? (-10'hc) : (15'h16)), w2, ((28'ha) ? w48 : (8'h1b)), $signed(w62), $unsigned(w60), (w83 ? w95 : w82), (!w73), (^(10'h8)), {w67, w93, (-27'h14), w99, (22'hf), w67, (-10'h6), w60, w42, (-29'h9), w68, w58, (-12'h1c)}} ? (|((^~(12'h4)) ? {(-27'hf), w62, (-2'hb), (21'h7), w5, (5'hb), w72, w51, (-18'h1), w64, w55, w3, w64, w98, (30'h13), (-25'h1a), w6} : (~|w68))) : {((-8'he) === w86), (+w85), (^~w61), $signed(w94), ((29'h19) ? (24'h11) : (27'h17)), $signed(w55), ((-8'hc) ? w75 : (-24'he))});
assign w41 = w5;
assign w42 = (~|((-w83) ? $signed((w90 ? (-22'h16) : (4'h3))) : (-26'h1b)));
assign w43 = (w45 << (-24'h15));
assign w44 = $unsigned(($unsigned($unsigned({(33'ha), (-25'h18), w85, (11'hb), w53, (32'h7), w64, (-10'h5), w62, (24'h3), w46, (8'h8), (8'hd)})) ? {w84, (14'h1b), (25'h1b), w93, (14'h5), (2'h1c), w49, w5, w1, (13'h1d), w57, w57, (-16'h6), (30'h1b), (9'ha), w52, w61, (3'h9), w85, (25'h1c), w71, w75, w49} : (18'h1e)));
assign w45 = (1'h8);
assign w46 = ({(+(2'h10)), {(7'h6), (-1'h5), w96, w78, w10, w62, (-22'hf), (-5'h8), (-17'h7), w90, w67}, (~^w98), (15'h2), ((10'hb) | (-21'hc)), (w74 ? w81 : w84), $unsigned((-4'h14)), {(-7'h3), w77, (-20'h13), w82, (-7'h8), w97, w60, (30'ha), w87, (-5'h11), w48, w81}, ((-7'h14) >> w10), ((28'h1d) ^ w100), {(-2'h1d), w76, (7'h16), w100, w93, (-15'h7), w94, w98, (-24'h12), w3, w90}, w73, w94, $signed((-24'hb)), w73, ((30'h1b) ^ (24'h11)), $signed((-8'h1c)), (29'h15), $unsigned((-15'h16)), (w61 ? w47 : (19'hd)), ((3'h1a) ? (-21'h13) : (7'hd)), (w68 === w83), w2, {(4'h16), w58, w89, w67, w80, (-11'h1e), w67, (-19'h12), (25'ha), (2'h18)}, (3'h8), (!w7), $signed(w2)} ^ {(27'h16), ((6'h19) ? (6'h4) : w92), ((-1'h13) ? w7 : w99), {w95, w58, w59, w95, w95}, w98, w98, {w87, (-22'h19), w10, (-14'h6), (3'h11), (-6'h1d), w52, w57, w48, (-20'h13), w83, (-5'h18), (-4'hb), (6'h1e), w7, w97, w100, w64, w58, w51, w97, w99}, (^~w65), w58, (~&(-5'h11)), (-10'h16), (~^w88)});
assign w47 = ((((w62 ? (17'h17) : w1) ? w8 : {(3'h2), (-12'h1), w94, (14'h14), (3'hb), w86, (14'h8), w83, w65, (-23'h4), w83, w49, w5, (7'h10), w77, (-29'h6), (-27'h1e), (-18'h18), w53, (-17'hd), w5, (-30'ha), w99, w66}) ? {(-30'hc), (-17'h9), w91, w50} : (-23'h0)) ? $unsigned(w52) : (12'h19));
assign w48 = (-18'h18);
assign w49 = w79;
assign w50 = ((^(w57 ? w53 : (18'h8))) ? (^w64) : (-15'h2));
assign w51 = (-7'h4);
assign w52 = {(~|(~^(28'h1c))), $unsigned({(-10'hb), (-2'hf), w57, (7'h6), w57, w89, w72, w61, w56})};
assign w53 = w96;
assign w54 = w85;
assign w55 = {(15'hc), (|(-16'h11)), {(33'h2), (-17'ha), (13'h14), (18'h3), (-25'h18), w7, (-2'h8), (11'hd), w81, w82, (-17'hb), (18'hd), w65, (-6'h17), (-21'h3), w99, w75, (-10'h1d), (21'h19), w77, (2'h2), w9, (-6'h18), (-20'h3), (-20'h18), (28'hd)}, $unsigned((^w62)), {w6}};
assign w56 = (w89 ? (!(~^(~|(w4 << w5)))) : ((20'h6) ? $signed((-23'h7)) : w76));
assign w57 = ((((-19'h11) === w65) ? ($signed(w65) ~^ $unsigned((-3'ha))) : (w96 - w93)) ? ({(-1'h5), (2'h1b), (-5'h15), w68, (19'hb), (-27'h13), (11'h7), w91, (22'h8), (-23'h18), (-7'h9), w9} ? $signed((10'h3)) : (17'h16)) : $signed({w63, (-2'h19), w89, (20'h14), w2, (-28'h16), w7, w3}));
assign w58 = $unsigned({$unsigned(w76), (~|(-12'h12)), (23'ha), {w7, (-2'h12), (-1'h0), (8'h1a), (24'hc), (28'h5), w81, w7, (-3'h11), w71, w79, (-26'h11), w7, w76, w75, (27'h7), w4, (6'hd), w89, w3, (-12'h1a), w84, w95}, (w88 ? (25'h12) : w85), $unsigned((-4'h7)), (^(8'h1d)), (w65 << (-14'hb)), (w61 * w68), $unsigned(w98), (-(-28'h11)), w1, (-24'h9), ((-24'h6) | (-29'h1c)), ((10'h12) == w64), $signed((8'hb)), (17'h4), (w75 ? (-17'h19) : w62), w65, (24'h1d), {(-19'h14), (-15'h15), w64, (-4'h6), w8, w70, (-4'h15), w69, (25'h16), w65, (25'h1c), (12'h9), (-23'h18), w1, (30'h18), w5, w60, w69, w82, w67, w3, (17'h16), w78, (7'h4), (-17'h17), w87}, $signed(w80), (-13'h1c), (+w6), (-w82), (15'h5), (~^w80)});
assign w59 = w95;
assign w60 = (w68 ? $signed($unsigned((+(!w100)))) : {w84, (!w3), ((30'h13) * w4), {w7, (26'h12), w9, w77, w95, (-7'h4), w94, w91, (5'h5), w91, w75, (-10'h1a)}, (-24'h9), w99, (w85 ? w81 : (27'hb)), (w8 ? (18'h8) : (25'h5)), ((-5'h17) ? (-3'h1c) : w10), w72, $unsigned((-2'h18)), {w3, w100, w69, (30'h8), w62, w96, w76, (20'h1c), w3, w99, (11'h1a), (-25'h3), w64, w74, w66, w94, w72, (9'h14), (26'h12), (-30'h18), (11'h19), w10, w86, w3, w63, (11'h11), w76, w97, (-25'hb), w80}, ((-15'h15) ~^ w64), $unsigned((-17'h8)), {w10, (-18'h9), (10'h13), w69, (21'h10), (1'h1e), w61, w72, w93, w67, (-8'h5), w66, (4'he), (18'hc), (20'h9), w79, (25'h14), (19'h4), w98, (-24'h2), (-20'h4), (-12'h5), (1'h7), (-18'h7), (8'hf), w8, w86, (-23'h1), w78, (-2'h1a)}, ((15'h10) ? w69 : (29'h11)), {(-15'h1b), w85, (19'h1), w5, w69, w69, (16'h1c), (-1'h15), (7'h12), (-9'h1b), (10'hf), (-6'h9), (5'h1e), w90, w84, w73, w91, (15'h9), w65, w74, (18'h2)}, (~|w66), $unsigned((-20'h19)), (-14'h9), {w71, w81}, ((17'h19) * w70), w91, ((-22'h11) ? (14'h3) : w79), (w93 ? (14'h15) : (-15'h8)), ((-31'h7) ? w1 : w75), (16'h13)});
assign w61 = (13'hd);
assign w62 = (~|(^{w65, (-18'h1e)}));
assign w63 = (~^w73);
assign w64 = ({(+w65), $unsigned(w73), (-(19'h1b)), (!w75), $unsigned(w100), (w84 >= w69), $unsigned((-2'h1b)), ((-17'ha) + (-15'h0)), (-20'h11), (-13'h13)} ? (w75 << $unsigned((-28'h7))) : ((-26'hd) ? w69 : w2));
assign w65 = {w89, (|w86), (^~$unsigned((29'ha))), ((w7 < (5'hd)) ? {w93, (20'hb), w81, w93, (19'h1d), (-18'h10), w8, (-27'h1b), w2, w79, (5'h5), w67, (14'h1a), w93, w81, w73, (-20'h1d), (16'h2), (1'h7), w87, (6'hb), (17'h18), (-27'hc), w75} : {w82, w75, w85, w5, (-20'h9), (-9'h18), w3, w93, (13'h18), (12'hc), w74, (-6'h5), (-1'h1c), (-26'h5), w91, w80, w95, (-25'h1c), (-24'h0), (8'hb), w95, (4'ha), w82, (-13'h9), w83, w6, (-3'h5), (15'he)}), $signed((|(-22'h5)))};
assign w66 = w67;
assign w67 = {{w70, (-3'hb), (5'hd), (28'he), (31'hd), w70, w93}, $unsigned((~^w96)), ((w7 ? (-10'h1a) : w80) ? ((21'hd) ? (-31'h1b) : w82) : $signed(w9)), (((-20'h17) ? (26'h1b) : w69) - (w4 ? w84 : w98)), $unsigned(w6), $signed(((5'h1b) ? w5 : w84)), (22'h11), {(24'h3), (-30'h1e), w79, w10}, $unsigned((w71 | w10)), (7'he), (-{w10, (-15'h14), (-8'h11), w82, (16'he), (2'h5)}), $signed((-4'h16)), (~&((4'h14) <<< w93)), {(32'hb), w79, (20'h16), w80, (18'hd), w78, w71, w96, (-23'h19), (-23'h16)}};
assign w68 = w9;
assign w69 = ((w83 | ((26'h7) ? (30'h4) : ((-6'h14) >> w1))) ? $signed(w1) : $unsigned((~|(|{w77, w72, (3'h3), w80, (7'h15), (-8'he), w78, (-13'h1)}))));
assign w70 = $signed(w88);
assign w71 = (|{$signed((-26'h10)), ((17'h18) ? w94 : w85), ((-29'h4) ? (-12'h9) : w89), (w8 ? w80 : (31'h15)), $unsigned((-9'h9)), {w89, w88, (-31'h1), (32'h15), w79}});
assign w72 = $signed((^{(-21'h11), w96, (-32'h13), (-6'h9), (12'h6), (17'h1e), w4, w86, (-8'h3), (-27'h16)}));
assign w73 = {{w84, (2'h9), w90, w1, w86, (-18'h17), w78, w90, (20'h15), w84, w94, (-3'h1c), w83, (7'h3)}, $unsigned((16'h1a)), ((|w9) ? ((8'h6) < w83) : (-25'h3)), {(7'h10), (-24'he)}, w3, ($unsigned(w92) > (27'h15)), w96, $unsigned((^w1)), w4, {(5'hf), (-5'h5), w4, w97, w84, w88}, (-9'h1d), {w85, (15'h1e), w9, (-20'h1a), w82, w99, (-15'he), (24'h11), w99, (29'h6), (13'h18), w6, (9'h1e), (-1'h16), (13'hc), w87, (-1'he), (-22'h1)}, {w8, (28'h1a), w95, (12'h12), w8, w95, w3, (-25'h1b), w84, w8, (25'hb), (-25'h9), w95, w83, (-19'h1a)}, ((!(-26'h1d)) ? {w88, (18'h10), (-4'h1d), (30'h4), w96, (18'h17), w100, w83, (27'hc), w7, w89, w85} : {(10'h12), (-15'hc), w90, w100, w99, w100, (-28'hc), (17'h1), (18'h3), w83, (-2'hc), (3'h7), (5'h6), w3, (30'h1a), (28'hc), (12'h8), (-7'h2), (6'h17), w1, w92}), {w85, (-29'h19), (30'h15), (5'h11), w10, w1, (-23'h7), w82, w98, w100, (18'h1), w10, (24'h1c), w7, w92, w95, w8, (2'h17), (33'hc), w9, (7'h1b), w7, w80}, (|((-2'h11) ? (13'h6) : (-2'h1b))), w97, (((9'h1) ? (-28'hc) : w85) ? (|(-4'hd)) : $signed((28'hd))), (-10'h1b), {(-17'h8), w6, (-23'h4), (16'hb), w96, (17'h12), w89, (-19'he), w83, (-14'h0), (-31'hb), (2'h13), (-31'hf), w3, (-32'h1d), (-21'ha), (12'h12), w96, (-24'h7), (15'ha), w83, (9'he), w80, w4, w84, w6}, (((-4'h10) ? (26'h3) : w76) ? (~^w80) : (!w77)), (-3'h3), w4, $signed($unsigned(w95)), ($unsigned(w4) == (-27'h7)), ((-(-14'h13)) ? (10'h9) : (w7 ? (33'h12) : (27'h3))), (((-15'h12) ? (-25'hd) : (26'h6)) != (^w84)), ((w77 ? (-27'hd) : w7) ~^ w89), (~^$unsigned(w79)), ($unsigned(w80) >>> (w6 ? (-10'h7) : w82))};
assign w74 = $signed({(|w88), {(-6'he), (-6'ha), w91}});
assign w75 = w8;
assign w76 = (-24'hb);
assign w77 = ((~|(20'h14)) ? w87 : (~&(&(+((-25'hb) && w9)))));
assign w78 = w89;
assign w79 = $signed(w87);
assign w80 = (w85 ? $signed({(-23'h10), w96, (6'h12), w89, (-3'h18), w97, w87, (26'hc), w92, w98, (-5'h1b), (-15'hf), w90, (12'h2), w96, w84, (22'h16), w1, w1, (27'ha)}) : (28'h5));
assign w81 = {$unsigned({(-22'h8), w8, w3, (-18'h8), (-28'h5), w83, w90, (-17'h1d), w1, (-28'h5), (-25'h19), (-27'h2), (-25'h11), (-19'h3)}), (-8'h11), {w88, w4, w3, (-2'hd), (11'h15), w100, w95, w90, (-2'hb), (28'h8), (-30'h0), (1'h19), w5, (-5'h5), w86, (5'h7), (-9'h13)}, ($unsigned((-13'h12)) != (-17'h19)), {w9, w93, w10, w100, w90, w10, (-26'h14), (8'h7), (-5'h1b), w84, w1, w92, (13'h18), (22'hf), (-18'h1), (30'h10), (23'h5), w93}, $signed($signed((-24'ha))), (~^(-w96)), (-23'h1e), ((-26'h12) + $signed((21'he))), w82, (&(-11'hc)), (!(+w90)), {w91, w89, w90, w94, (3'h1a)}, {(-27'h14), w89, w5, (12'h18), (19'h10), (-9'h19), (19'h3), w91, (-3'h6), (-9'h13), w4, w93, w99, (25'h2), w94, (-27'ha), w8, (-19'h18), w8, (19'h2), w91, w98, w94}, $signed(w7), w1, (!((11'hf) ^ w10)), (13'h1d), {w1, (-15'h11), (34'h11), (19'h14), w82, w94, (16'h8), w92, w3, (-22'h6), (-28'he), (-11'h17), w92, (9'h8), w90, w100}, (!{w82, w2, (5'h14), w4, (20'h8), (-9'h19), (30'h17), w82, (9'h1b), w8, w3, w4, w98, (-27'hd), w9, w96, w89, w88, w91, (-8'h13), (-32'h1), (-30'h8), (-24'h5), w98, w7, w85, w87, (-33'h4)}), (~&$signed(w6)), (19'h4), (!(^~w90)), w8, {(10'h13), (-10'he), w99, (-16'h5), (-12'h17), (-12'h1a)}, w83, (-29'hf), {w10, w83, w87, w82, w4, (30'hc), (-3'ha), w1}, (-4'h1a), ((w4 + (8'hb)) <<< ((-10'h0) ? (11'h12) : (14'h7)))};
assign w82 = (~&{{(-27'he), w93, w3, w86, w10, (-20'h14), w98, (4'h1), (18'h12), w98, (6'h1c), (-22'h12), w87, w4, (6'hd), w84, w10, w83, (-37'h16)}, w92, (w88 ? (29'h1) : w83), (+w93), $signed(w97), {(-22'h12), w84, w97, (-22'h15), (24'h1e)}, ((-30'h1c) >> (-1'h17)), (w93 ? w6 : w88), w90, $signed((11'h3)), ((26'h2) ? (-13'h8) : (-4'h1c)), w86, (w97 ~^ (-3'h17)), (9'h3), {w86, w87, w6, w92, w98, (29'h1d), w88, w4, w96, (-23'h6), (10'h14), w100, (15'hd), (8'h5), w100, w2, (3'h19), (-8'h6), w4, w96}, (7'h19), $signed((16'h1d))});
assign w83 = (1'h1c);
assign w84 = ((-18'h1d) ? (~&(((-3'h9) ? (-28'hf) : (25'h1d)) ? w93 : (4'h1))) : (+((~|{w91, w97, w6, (-16'h1b), (21'he), w91, (-12'hd), (-31'h9), (8'hc), (-15'h8), w8, (-31'h15), w98, w92, (-28'h1e)}) ^~ {w90, w2, w97, (-14'h9), w2, w98, w90, w95, w99, w7, (14'h12), w8})));
assign w85 = (-21'h19);
assign w86 = ({w5, w90, {w9, (-27'h8), w93, (-14'h1d), (-20'hb), w10, (-5'h17), w91, w10, (-25'h1c), w100, (32'h1c), (27'h12), w99, w93, (4'h5), w99, w87, w4, (-22'h18), w93, (-24'h1c), w91}, ((-4'h1a) && w94), $signed((-2'h1)), ((6'h4) ? (22'hd) : w94), {w98, (26'h1), (16'h2), (31'h13), w100, w98, (-28'hd), (19'h17), (-5'hc), (-25'h1d), (13'hb), (-18'h14), (12'hb), w88, (-11'h10), w2, w97}, (30'h14), {w10, w4, (19'h7), w97, w6, (27'h1), (21'ha)}, (!w6), ((-5'h1d) >> (-28'hc)), (-1'h6), $signed((4'h7)), (w98 != w91), (-31'h6), {w9, (-20'h2), (-17'h13), (7'h12), (20'h1), w94, w1, w93, w93, w97, (5'h7), w94, w4, w94, w3, (-8'hc), w9, w100}, {(3'h1d), w9, (30'hf), (-30'h14), w92, w100, w90, (-3'h18), w5, w98, w97, w8, (9'h1e), (-20'h4), (11'h12), (29'h7), w89, w96}, ((18'hf) ? w5 : w5), (w7 | w88), $unsigned((23'h19)), (^~(-8'h1b)), (w92 ? w87 : w8), {w4, w100, w97, (28'h15), w89, (-29'h1), w92}, (w89 ? w5 : (8'h1b))} ? {$signed(w95), ((15'h1c) ? w9 : (7'hd)), $unsigned((32'h5)), ((29'h16) ? (30'ha) : w90), {w98, w9, w95, (-10'he), w90, w6, w93, w1, w3, w8, (9'h6), (-25'h6), (12'h18), (3'h4), (-5'hb), w89, w4, w4}, $unsigned((15'h11)), (w7 ^ w97), (30'h14), ((6'h2) ? w98 : w91), (-w92), (w3 ? w90 : w2), ((12'h19) === (-14'hf)), {w93, w88, (20'he), w93, (-16'h4), w100, w6, (-2'h2), (5'hf), (26'h1b), w6, (12'h16), w6, (-11'h5), w7, w87, w89, (23'h2), (5'h1d), (-12'h9), w4, (-30'h1e), (10'hf), w92, (-5'h16), (-14'h3), w88, (-6'ha), w96}, ((19'h9) ? w92 : w6), (^w94), ((19'hc) ? w97 : (27'h3)), (18'h14), (~&w93), {(9'hd), w3}, $signed(w3), (-13'h5), (w97 + (-2'h6)), (^w6), (29'h10), {(-22'h6), (-15'h8), (21'h16), w9, w2, w97}, w95, $unsigned((-15'h3)), (20'ha), ((-21'h1c) ? w88 : (-14'hf))} : w3);
assign w87 = $signed((w88 << (-22'h2)));
assign w88 = (!{((-26'hd) ? (-5'hb) : w5), ((24'h1d) ~^ (16'h15)), (&(21'h9)), ((-12'h11) <= (-5'h14)), (w89 ? (-20'h4) : w96), (&w5), w10, (~&w4), w92, {w91, (-29'h1a)}, (&w7), ((18'h15) ? (17'h8) : w93), (^(29'h1e)), {(16'h17), (-32'h12), w7, w10, w91, (13'he), w4, w6, w96, (9'h1c), w1, w1, (-25'h17), (17'h9), (-24'h4), w1, w7, w94, (20'h19), (-4'h1), w99, (-22'h7), w100, (-19'h1a), w8, (19'h1c), w97, w9, (-26'hc)}, ((-19'h11) ? (17'h8) : (-18'h2)), (-9'h16), $unsigned((-12'h1)), {w6, w1, (22'h11), w10, w99, w95, (23'h5), w100, (-15'h5), w100, (10'h1b), w90, (-5'h9), (-15'h1a), w5}, $signed((2'h15)), w100, (w90 - w98), (w3 & (23'ha))});
assign w89 = (^~(({(3'h18), w100, (-22'h18), w97, (1'h1e), (-1'h5), w100, (28'h3), w10, (14'h6), (11'h9), (-4'h8), w93, (-26'h15)} ~^ {(-18'h1), (11'h13), (10'h1a), (2'h3), (-36'h2), w91, (-17'h7), w9, (18'h4), w8}) === w100));
assign w90 = (w2 ? $unsigned($signed({w91, w97, (-20'h1a), (-17'h0), (-1'h1d), (-8'h5), w96, (1'h5), w100, (-21'h3), (10'h1e), (9'h11), w10, (-26'h12), (8'h2), (20'h6)})) : w7);
assign w91 = ((-21'h1a) ~^ w8);
assign w92 = $unsigned(w100);
assign w93 = w2;
assign w94 = {((^~(30'h16)) === (w7 ? w98 : (-17'h18))), w98, (!(~|(-16'h1a))), {(22'h4), (-18'h1), (-23'he), w96, w96, w8, w3, (28'h3), w10, (-15'h1), w7, (11'hc), (-27'h4), w5, w100}, (&(w100 ? (-18'h7) : (-30'h10))), (&(w100 - (12'h10))), {w4, (-32'h8), w96, w7, w3, w9, w5, (30'h4), (27'h14), w100, (-23'h9), w100, (-22'h12), w3, (6'hd), w9, (-27'h10), (-34'h1d), w98, (1'h19), w8, (34'h4), w4, (-6'h9)}, ((~|(-15'h11)) == (~&w98)), (((-25'h6) < (-30'h12)) ? (^~(-5'hb)) : (w8 ? w96 : (15'h2))), (+{w10, w99, w2}), ((19'h4) - (&w7)), w1, ((~^w7) ? ((4'h1b) ? (-19'h16) : (-5'h14)) : (w2 ? w2 : (-8'h13))), (w5 ? $unsigned((-8'h18)) : {(21'h3), w7, w3, (-10'h9), w95, w8, (-1'h14), (25'h2), (3'hf)}), (~|(-2'hb)), w99, (!(-23'h1c)), (22'hb), ((^~w96) ? (w95 ? w1 : w7) : w2), {(10'h4), (-5'h11), w96, (4'h7), w100, (17'h8), w97, w10, w97, (-14'h2), w7, (-26'h14), w2, (-7'h16), (8'h1e), (-7'hf), w5, w10, (1'h13), (9'h1), (19'h4)}, (((-7'h1a) ? (3'h1e) : w100) >>> $unsigned((29'h14))), w100, {w98, (-30'h16), (-21'h18), (-8'h3), (23'h14), w97, (2'h17), w98, (2'h10), (-1'h16), (16'h1e), (20'h1d), (16'hb), w100, w6, (-4'hc), w8, (25'hf), w4, w96, (23'h6), (22'h19), (-29'hc), w9, w5, w97, w97}, $signed((+(-11'h11))), (~^((31'h7) >= (22'h5))), ({(-9'hd), w99, w9, (-27'h2), (9'h14), (15'h12), w6, (11'h1), w98, w6, (-3'h13), (17'ha), w9, w5, w95, (29'h15), w10, (29'h2)} ? {(-20'h1a), (20'h1b), w1, w97, (-3'h15), w2, w8} : (-11'h3))};
assign w95 = ($signed(w5) << (14'hc));
assign w96 = (-2'ha);
assign w97 = (-9'hd);
assign w98 = ((-(5'ha)) ? {(w100 ? (3'h19) : (14'h12)), ((-14'h13) <<< w100), w99, (&w3), {(5'h5), (7'h16), (-24'hf), w99, w8, w4, (10'h1e), w4, w10, (-17'h1a), w3, (-9'h1c), (16'h1b), (29'hd), w8, w9, (17'h1b)}, $signed(w4), ((11'h15) & (32'h10)), (w3 ? (19'ha) : w8), w1, ((16'h15) !== (27'h1b)), ((21'h5) ? w6 : (-9'h1)), $unsigned((10'h1d)), w9, (w7 ? (-4'h17) : (-10'h2)), {w4, (23'h9), w8, (-27'hc), w1, (-28'h0), (21'h11), w99, w5, w2, (-5'h0), w1, (31'h1d), (-16'h11), (-19'h1c), w100, (-23'h19), (14'h1b), (-4'h6), w100, (7'hf), (-7'h10), (13'h17)}} : ({w9, (-22'h1e), w6, w8, (-14'hf), (26'hb), w1, (-19'h13), w4, w4, w1, w99, (-16'hd), w100, (6'h6)} ? w3 : (-19'h12)));
assign w99 = ({(17'h19), {w3, (5'h9), w4, (15'hc), (-30'h18), (-5'h14), (27'h15), (24'he), w10, w8, w2}, w4, w1, ((-18'h13) - (-25'h9)), (~|w2), ((8'h1e) ? (-17'hf) : (-13'h9)), (w7 >= (-13'h6)), (-23'hd), (4'h13), (w8 >> (-11'h14)), w3, w8, {(-4'ha), w8, w10, (21'h1e), w100, w5, (-18'h16), w100, (7'h6), (12'h5), (14'h13), (-26'h7)}, (w6 ? w6 : (-13'h13)), (w5 ? w10 : w100), w2, w4, (4'h5), (11'h15)} ? $signed((|(17'h1e))) : $unsigned((~^((-7'he) ^ {w100, (-7'h10), (-13'h7), w9, w3, (-10'h13), (3'h17), w6, (21'h6), (-29'h6), (28'h19), w1, (-19'hf), w10, (7'h12), (26'h9), w7, w6, w100, (-21'h15), (18'hb), (-6'ha), (16'h16), (12'h17), (-6'h17), (-7'h15), w1}))));
assign w100 = (-10'h17);
assign y = {w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100};
endmodule
