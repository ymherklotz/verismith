module test_module(y, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10);
output wire [1372:0] y;
input wire [6:0] w1;
input wire [18:0] w2;
input wire [9:0] w3;
input wire [5:0] w4;
input wire w5;
input wire [28:0] w6;
input wire [17:0] w7;
input wire [29:0] w8;
input wire [10:0] w9;
input wire [5:0] w10;
wire [20:0] w97;
assign w97 = ({(w9 ^ w7), ((-(27'he)) != (1'h0)), ((-(19'h17)) ? w1 : (23'h1e)), (w10 ? w9 : (1'h11)), (w2 ? (1'hc) : (8'h5)), (-(28'h11)), (w3 ? (1'h0) : w6), $unsigned(w9), ((1'h0) > (-(5'hc))), (-(5'h14)), ((-(20'h0)) ^~ (-(4'h1b))), {(8'ha), (1'h0), w1, (-(3'h1d)), (1'h0), w6, w9, (-(15'hc)), (1'h0), (-(18'h4)), (-(4'h1b)), w3, (20'h6), (27'h5), w3}, (1'h0), (~^(-(26'h11)))} ? $signed(($signed((-(7'h1c))) ? (w4 >>> (-(2'h4))) : ((-(23'h10)) && w3))) : {(+(-(17'he))), (^(18'h10)), {w2, (1'h0), w7, (1'h0), (-(26'h1)), w6, w4, (9'hb), (29'h1), (-(1'h1e)), (-(15'h11)), (29'h18), (-(4'h1a)), (23'ha), (24'h14), (17'h10), (28'h14), (32'hc), (1'h0), (-(29'hc)), (-(10'hf)), (-(24'h11)), (31'h19), w2, (-(14'h15)), w6, w4, (2'hc), w7, (-(17'h7))}, (&(1'h0)), {(29'h18), (-(25'h4)), (6'h13), (27'h7), (-(22'h18)), (-(23'h4)), w3, (-(26'h1)), (29'h1d)}, ((19'h1b) ? w3 : w3), (4'ha), $unsigned(w6), ((-(19'hc)) ? w8 : (29'h9)), (1'h0), (w7 && w4), (|w5), {(7'h4), w1, w3, (1'h0)}, w10, ((-(2'h13)) * (1'h0)), (w8 + (-(5'h12))), (-(17'h16))});
assign y = {w97};
endmodule
