module test_module(y, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10);
output wire [1328:0] y;
input wire [19:0] w1;
input wire [5:0] w2;
input wire [29:0] w3;
input wire [20:0] w4;
input wire [7:0] w5;
input wire w6;
input wire [18:0] w7;
input wire [11:0] w8;
input wire [20:0] w9;
input wire [26:0] w10;
wire [11:0] w11;
wire w12;
wire [1:0] w13;
wire [16:0] w14;
wire [28:0] w15;
wire [28:0] w16;
wire [16:0] w17;
wire [1:0] w18;
wire w19;
wire [4:0] w20;
wire [26:0] w21;
wire [25:0] w22;
wire [11:0] w23;
wire [9:0] w24;
wire [7:0] w25;
wire [22:0] w26;
wire w27;
wire [25:0] w28;
wire [16:0] w29;
wire [8:0] w30;
wire [29:0] w31;
wire [17:0] w32;
wire [11:0] w33;
wire [16:0] w34;
wire [7:0] w35;
wire w36;
wire [9:0] w37;
wire [22:0] w38;
wire [1:0] w39;
wire [9:0] w40;
wire [21:0] w41;
wire [29:0] w42;
wire [20:0] w43;
wire [3:0] w44;
wire [16:0] w45;
wire [21:0] w46;
wire [20:0] w47;
wire [6:0] w48;
wire [4:0] w49;
wire [2:0] w50;
wire w51;
wire [8:0] w52;
wire [5:0] w53;
wire [18:0] w54;
wire [14:0] w55;
wire [14:0] w56;
wire [26:0] w57;
wire [9:0] w58;
wire [6:0] w59;
wire [27:0] w60;
wire [13:0] w61;
wire [11:0] w62;
wire [17:0] w63;
wire [15:0] w64;
wire [24:0] w65;
wire [6:0] w66;
wire [8:0] w67;
wire [27:0] w68;
wire [13:0] w69;
wire [15:0] w70;
wire [4:0] w71;
wire [25:0] w72;
wire [2:0] w73;
wire [17:0] w74;
wire [16:0] w75;
wire [22:0] w76;
wire [11:0] w77;
wire w78;
wire [18:0] w79;
wire [10:0] w80;
wire [22:0] w81;
wire [26:0] w82;
wire [25:0] w83;
wire [16:0] w84;
wire [8:0] w85;
wire [25:0] w86;
wire [20:0] w87;
wire [18:0] w88;
wire [17:0] w89;
wire [9:0] w90;
wire [22:0] w91;
wire [26:0] w92;
wire [11:0] w93;
wire [19:0] w94;
wire [2:0] w95;
wire [25:0] w96;
wire [14:0] w97;
wire [6:0] w98;
wire [10:0] w99;
wire [1:0] w100;
assign w11 = $unsigned($unsigned((+({(-16'h1a), w23, w89, (25'h14), (4'h19)} ? ((-18'h16) - (-26'h12)) : $unsigned(w43)))));
assign w12 = ({(w47 >> w43), w68, ((20'h10) ? (-23'h1b) : w27), (w83 ? w7 : (21'h17)), (+w54), {(22'h5), (5'he), (22'h1a), (27'h2), w18, w54, w69, (-28'hb), (-28'he), w92, (16'h3), (-4'h1d), w47, w13, w82, w43, w83, w37, w10, (14'hc), w64, (11'h3), w45, w54, (-4'h8), w76, (30'h9)}, w58, (-11'h1b), w9, w61, {w18, (20'h17), w78, w77, (16'h1b), (25'hb), (13'h19), (19'h17), w24, w38, (25'h15), w40, w66}, w3, (w32 <= w91), w64, ((10'h1e) ? (7'h4) : w99), ((19'hf) ? (-13'hf) : w36), (w90 + w22), (~|(12'h19)), (w61 <= w40), (w49 ? w50 : (23'h6)), ((-12'ha) ? w33 : w3), ((-20'h5) ? (-22'he) : (26'h10)), (!w59)} ? (({(-5'ha), (-20'h1a)} - w44) + (!$signed($signed((-33'h12))))) : (w40 ? (w3 ? w69 : ((-1'h5) ? w24 : (-18'h12))) : $signed($unsigned(w9))));
assign w13 = (|w28);
assign w14 = (-19'hf);
assign w15 = {((24'h19) || (^~w34)), {w50, w49, w99, (15'h3), (-7'h3), w7}, ((-20'h6) >>> ((-16'h1e) ? (-11'h16) : w60)), $unsigned((~^(2'h7))), w66, ((w77 ? w5 : (-5'h4)) ? (-6'h15) : {(20'h1d), (-25'h2), w90, (16'hd), (22'h10), w36, (-20'h14), w77, (-24'hb), w74, (-7'h10), w10, (1'h1e), (20'h7), w50, w5, w3, (-17'h12), w38, (18'hb), (32'h11), w90, (21'h11), (-5'h8), w84, w44}), {w92, w47, (7'h3), (-29'he), (23'h1d), w51, (-19'h17), (-26'h5), (25'h2), (-32'h13), (-26'h1a), w85, (-26'h14), (21'hf), w5, w55}, (-22'h16), (~^(w3 >= (32'h1e))), w38, (-7'h19), (30'h12), w16, ({(-24'h14), w41, w74, w78, (19'h2), w35, w18, (28'h6), w90, (-24'h10), w51, (-6'h1a), (-14'h19), w92, (-9'h3), w66, w43, (11'h3), (27'hf), w98, (6'h5), w71, w42, (9'ha), (-23'hd), w87} <= (+(-25'ha))), ($signed((19'h3)) ~^ (-w7)), (~&w56), {w95, (-24'h1c), (-2'h1), (25'h1e), w72}, $signed((w93 << (-11'h16))), w19, {(-28'h3), (29'h1), w54, (5'ha), (1'he), (4'h1c), w89, (-30'h2), w56, w74, (3'h16), (-18'h16), w30, w19, (27'h1d), w9}};
assign w16 = {w71, ({(-25'h16), w64, w66, w95, (16'h6), (18'h9), w6, (-16'h1c), (-16'h1a), w6} <= (10'h14)), w27};
assign w17 = w83;
assign w18 = w30;
assign w19 = ($signed((^((26'h1e) ? (~&w61) : (5'hf)))) >> (^~w92));
assign w20 = w81;
assign w21 = (-15'h1d);
assign w22 = {(7'h13), {w33, (-14'h1c), w9, w45, w59, w51, w68, w51, (-17'h10), w86, w35, (-11'hb), w36, (17'hb), (14'h13), (-5'hb), (11'h8), w81, w71, w3, (-24'h12), (-30'h5), (-23'h5)}, (-25'h5), (|((19'h3) >= w59)), {(6'he), (-14'h13), w69, (-6'h1b), w86, (-20'h14), (-18'h11), w80, (-28'h6), w9, w68, (-12'h1e), (12'hb)}};
assign w23 = $unsigned((({w5, (-3'ha), w64, w49, (-6'h5), w30, (27'h1e), w39, w91, (6'h1d), w82, (16'h12), w38, w24, (-5'h2), (5'h13)} >>> ((-7'h3) ? w40 : w5)) ? $unsigned((17'h18)) : {w34, w34, w49, w90, (-6'h2), (-10'h19), (-29'h16), w33, (-16'h7), w52, (2'h3), (19'h13), (5'h2), (24'h3), w2, (-27'h1a), w77, w100}));
assign w24 = w58;
assign w25 = $signed($unsigned((3'hb)));
assign w26 = $signed((&((^~(w31 & (-10'h8))) ^ (!((8'h14) ? w35 : w55)))));
assign w27 = (23'h12);
assign w28 = ({$signed((17'h4)), w65, ((-20'h14) && w73), $unsigned(w4), (+w63), (15'h8), {w32, (16'h3), w95, w8, w68, (21'h5), w3, w90, (-23'h7), w41, (13'h1c), (-4'h2), (-17'h17), (-25'h17), (21'hc), (10'h5), (-25'h7), (-11'hd), (-1'h11), w32}, (w85 ^~ (21'h1b)), (w78 ? (28'hb) : (27'h14))} ? {((15'hf) ? (-28'h12) : w90), w63, {(21'hb), (19'h14), w40, (-21'h1d), w98, w10, w85, w54, w75, w81, w5, w8, (26'h19), w92, (10'h1c), (27'h1e), w83, w5}, w5, ((26'h3) >= (-28'h12)), (&w78), (|w58), w36, (-w84), w74, w98, (-13'h6), $signed(w37), $signed(w79), {w35, w76, w56, w34, w1, (-1'h7), (-6'h1d), (27'h9), (-22'h10), w8, w98, (-14'h15), (-24'h1d), (-13'h1c), (-3'h5), (-5'h3), (6'h2), (13'he), (17'hd), w35}, w89, w36, (|w77), w91, ((-26'h1e) ? (-9'hb) : w77), w93, $unsigned(w5), (~^w3), (+w68), (19'hc), (|w29), (-22'h1e), w80, $signed(w10), {w52, (-7'hb), w55, w73, w32, w30, (-32'h1c)}} : {((-9'h12) | (11'h17)), w86, {(-24'h1), (19'h5), w80, w82, (-11'h19), (7'h8), w42}, (w45 == (14'h17)), (-4'h6), $signed((21'hf)), $signed((-22'h18)), (-8'h12), (w58 >>> (-9'hb)), $signed((-4'hc)), w10, {w66, (5'h17), (-6'h2), (18'h9), (13'h2), (-11'h5), (-23'h1b), (-13'h4), w50, (-14'hb), w34, w90, w87, w71, w70, (-16'h1), (-6'h1e), (3'hd), (14'ha), w78, w66, (16'h17), w99, (7'h15), (6'h12), (-2'h4), (17'h19)}, (~&(32'h18)), (1'hb), $unsigned(w65), (w42 ? w62 : w55), w64, (29'h8), w73, {w45, w38, (2'h1a), w75, (-7'h10), (22'h9), (1'he), (23'h1e), (4'hf), (13'h12), w4, w71, w55, (30'h17), w74, (3'h11), (-17'h0), w76, (6'h1c), (14'h1), w4, (-11'ha), w84, w8, w32, (-29'ha)}, (4'h16), (+w99)});
assign w29 = $unsigned({(-15'h1d), (w85 !== w67), (w35 <= (11'h4)), ((2'h8) ? (19'h7) : (-27'h18)), (^~(22'h1c)), (~&(-20'h1a)), (18'h4), (w76 !== w54), w7});
assign w30 = $signed({{(26'h18), (17'h1), w94, w45, w56, (-25'h1c), (4'h12), (6'h12), (-1'h17), (4'h9), w3, (5'h5), (-1'h15), w54, w41, (23'h1b)}, (w62 ? (-13'h2) : (-22'hf)), {(-20'h8), w68, w1, w94, w80, (-10'h1b), (-5'h8), (19'hf), (-14'h0), (17'h1e), w99, (-11'h5), (10'h1e), w100, (-17'hb), (-29'h3), w97, (-29'h18)}, {w34, (1'h1c)}, w41, (w79 ? w95 : (-24'h11)), w43, (+(-12'h1d)), {(13'h1d), w43, w100, w83, (11'hf), (-4'hf), w99, (16'h1c), (-29'ha), w63, w75}, ((31'h19) == w95), ((4'h10) + (-28'h12)), w42, (w82 * w89), $signed(w94), {(24'hc), (-33'h15), w44, (-25'ha), (8'h13), w3, w31, (28'ha), w95, w68, w93, (-7'h13), (23'hc), w79, (30'h13), (-31'hc), w83, (18'h1d), w98, w54, w59, w49, w7, w61, w10, (-11'hf), (12'h10), (-14'h1), w62}, (w85 ? w35 : (24'h15)), (w4 - (23'h11)), (~|w37), (w90 ? w40 : (24'h10)), (~^(30'h4)), (w67 == w74), w80, $unsigned((-24'h4)), $signed(w55), {w7, (21'h1b), (6'h16), w50, (16'h14), (-25'h9), (-28'h12), w62, (-20'h15), w35, (24'h12), (9'h9), w100, (-11'h7), w4, w46, (-1'hc), (5'hd), (-11'h16), w98, w1, (-1'hb), w31, (-12'h7), (-5'hc), w1, (29'h13), w69, (-1'h7)}});
assign w31 = (^~(&$signed(($signed((-15'h13)) ? (~&(-25'h1)) : (w39 ? w50 : w35)))));
assign w32 = $unsigned($unsigned(($unsigned($signed(w6)) >= (13'hc))));
assign w33 = $signed(((+((w44 >> w98) === (w3 ? (2'h1) : (-34'hd)))) == {(25'h1c), w61}));
assign w34 = ((($unsigned(((3'h11) ? w69 : w93)) <<< {(-19'ha), (-23'hc), (25'h16), w2, w6, w51, w80, (-29'h16), (-14'h4), w53, w95, w66, (-32'h0), (-14'h1c), (20'h7), w78, (-12'h1c)}) ? $signed((^{w78, (-19'h8), (7'h2), (-20'h1d), w7, w59, (-12'h2), w82, (-16'h8), (15'h12)})) : $signed(((-8'h14) <<< w54))) == (|(+$signed((w98 >> w39)))));
assign w35 = (~&($unsigned(w74) ? $signed(w99) : {(4'h4), w78, w56, w3, w73, w82, (18'hf), w59, w59, w41, (27'h6), (-20'h1b), w78, (-25'h16), w10, (20'h14), w1, (-15'h3), w96, w64, w1, w44, w75, (3'ha), (-4'h11), w52, w83}));
assign w36 = w60;
assign w37 = (^{w61, {(-11'h1), (5'h19), (17'h8), (-19'h3), w75, (18'h2), (-10'h19), (-7'h1d), w48, w71, (-5'hc), (-10'h3), (-2'h16), w90, w10, w69, w89, w58, w62, w90, w3, w3}, w2, $unsigned(w85), ((-19'h1e) ? (-28'h18) : w67), {w84, (15'h1b), w4, w38, w4, w72, (-24'he), (-4'h0), (15'hd), w60, w100, (-20'ha), (-24'h7), w65, w95, w81, w97, (-21'h6), w56, (-22'h1e), (23'h11), (13'h1e), (15'h7), (29'h6), (-12'h1e), (-30'h1c), (11'h7), (5'h6)}, w73, $signed((-14'ha)), {(-26'h10), w46, (-17'hd), (18'h16), w92, (-25'ha), w82, (9'ha), w41, w4, w93, (29'h1), (9'h7), (-2'he), w80, w79, w85}, (!w61), (+(-2'h0)), {(22'h12), w58, w71, (-14'h6), (-11'he), w88, (-13'h1d), (-27'h19), w55, w38, w87, (23'h3), w71, w5, (27'h5), (-22'h1b)}, $signed(w61), ((-13'h3) - w91), (w73 ? (9'h4) : (26'h18)), (w94 ? w49 : (-10'hc)), ((-14'h5) ? w56 : (4'h18)), $signed((-31'h17)), (w7 ? w68 : (-28'h4)), $unsigned(w4), (-23'h4), (w44 ? w97 : (9'h12)), (-16'h1e), (w38 ? (8'h8) : (-8'h17))});
assign w38 = ($signed((-12'h13)) || $signed({w49, (-3'hc), w63, (-12'h14), (-29'h9), (18'hf), (-10'h16), w92, (-21'hc), w75, w42, w100, (-3'h1e), (-4'h9), (-5'h8), (-27'ha), (19'h1a), (18'h11), (-14'h14), (9'h1a), w97, (25'h4), w95, (9'hf), w7}));
assign w39 = {((21'h15) ? w57 : (12'h1)), w82, (-(&w72)), (-23'h9)};
assign w40 = w4;
assign w41 = ((~^{(24'h1), w57, w84, w6, (29'ha), (-8'h6), (19'h8), w2, (23'hd), (-14'h11), (17'h9), w80, (-20'h6), (-13'h1c), w94, (26'h1d), (31'h1c), (17'hf), (-29'h17), (-9'h1e), (-22'h1c), (31'h3), w69, w86, w92}) <= (4'h1b));
assign w42 = w2;
assign w43 = ((+(($signed((-15'h1)) ? ((18'h1b) << w46) : w86) !== $signed((~&(-2'h19))))) | (~&(w83 !== $unsigned((-20'h12)))));
assign w44 = {(!(3'h14)), $unsigned({w54, (5'h11), w94, (18'h3), w9, w98, (3'h7), (-8'h4), (-29'he), (11'h1), (12'h12), w74, (-2'h19), w46, w4, (-3'hc), (-21'h19), w48, w58, (-28'h9), (16'hc), w62, w53, (-25'h2), w61, w72, (-19'h1e), w46, (26'h1e)}), w84, $signed((+(7'h10))), (((-10'h1a) ~^ (-26'hc)) - {w52, (-17'h1a), w59, w96, (-28'h7), (27'h2), (31'h7), w56, (-7'h8), (1'h3), w88, w53, w76, (23'h16), w82, w62, w48, (-7'h1b), w50, (17'h15), (15'h15), (9'h10), (25'h15), w71, (-18'h16), (-29'h5), (10'h3), w77, w57}), (w62 ? ((-2'h1d) | (3'h7)) : w3), {(13'h11), w72, w77, (2'h1d), w87, (2'h16), w75, w89}, {(28'hb), w97, (-26'h0), w94, w87, (-16'h8), w60, (-12'hc), (3'h18), w91, (-20'h11), w99, w7, (24'h4), (-7'hb), (1'h15), (-30'h0), (16'ha), (-7'h10), w79, w45}, {(-21'hf), (-24'h13), (10'h19), w9, (11'ha), (-15'h1a), (-12'h1c), w83, (29'h8), w87, (-8'h13), (4'h4), w51, w64, (-5'h7), (4'h17), w85, w56, (19'h15), w4, (14'he), w8, w88, w75, w79, w82, (-19'h8), (11'h15), (-14'hb), (7'h19)}, (5'hc), (^(w82 ? (-20'h0) : (2'h6))), ({(-4'ha), (30'h1b), (-18'h1d), (-20'h19), (-9'h16), (-3'h1e), (-23'h15), w75, w85, (-24'he), w96, w46, w98, (-6'h11), (29'h2), (25'ha), (-24'h18), w73, w10, w48, w6, w1, (-1'h11), w81, w94, w79, w10} | ((-24'h1e) ? (-15'h1c) : (-16'h1e))), $unsigned((12'h1a)), w46, (+(&w83)), ((~|(-18'h17)) ? (w64 ? (-29'h3) : (-33'h1c)) : {(-29'h5), w99, (18'h8), (-18'h1), w79, w86, (-24'h13), w84, w8, (-5'hb), w92, w74, w92, w8, w2, w92, (-14'h19), w9, w47, w75, (4'h13), (8'h2), (-2'ha), w63}), (((-14'hd) ^ w75) ? (^~w75) : (w72 ? (14'h17) : w68)), ((w70 ~^ (-13'h14)) ? w66 : w46)};
assign w45 = {$signed(((8'h9) ? w56 : w63)), w98, {(-10'hc), (-27'h4), (-17'h1e), (-28'h1d), (-5'h12), w83, w68, (-21'hb), w55, w66, (-14'hc), (-21'h1e), (23'h2), w81}, {w95, (-24'h8), (29'ha), w80, (-7'h15), w71, w90, (-7'h9), (5'h17), w59, (-4'h1b), w98, w83, w98, (32'h3)}, (-18'h16), (~^(~^w10)), {w46, (5'h10), (8'he), w94, w100, w46, (29'h1c)}, ((~^w1) ? (|(-8'h1)) : (w81 ? (26'h18) : w9))};
assign w46 = w56;
assign w47 = $signed($signed($signed((~^$signed(w99)))));
assign w48 = (10'h7);
assign w49 = $unsigned({(9'h11), {(-23'h4), (-6'h8), w2, w84, w76, (-15'h1a), (27'h6), w8, (-6'h1c), w70, (-26'h1c), (-2'h15)}, $unsigned(w96), (-3'h1c), {(1'h19), w59, (-20'h2), (-1'h6), (-20'hb), w66, (30'h4), w1, (23'h1c)}, {w5, w8, (32'hb), (-9'hd), (4'h11), (-6'h0), (-31'h1a), (-29'hd), w65, w69, (25'hf), w71, w7, (2'hb), (22'h2), w74}, w71, ((19'h4) ~^ w55), w97, ((-24'h6) <<< (4'h1c)), (~^(-30'h17)), $signed(w82), {(12'h6), w57, (15'h19), (-18'h12), (-4'h3), w6, (20'h19), w86, (22'h14), (5'h14), w2, (29'h2), (-24'h10), w75, w71, w74, w89, w56}});
assign w50 = ((-9'he) ? (w94 < (26'ha)) : $unsigned(w59));
assign w51 = (7'h17);
assign w52 = {w92, $signed({(-6'h18), w67, (-25'hc), (23'hd), (-18'h19), w7, w65, (34'h1c), w5, (-5'h7)}), {(28'h1), (-8'he), (17'h1c), (-21'hb), (28'h3), (13'h8), (20'h8), (30'h8), w68, (-12'h10), (9'h1d), (-11'h7), w73, (-8'h7), w61, w97, w71, w98, w1, w78, w98, (29'h1c), (-27'h14), w94, w73, (7'h6), w95, (-24'h1d), (-17'hc)}, w79, w98};
assign w53 = ((&(12'h19)) | ({w57, w84, (29'h17), w80, w63, w93, (-31'h1d), w94, w9, (24'h2), w74} > (~&$signed((11'h2)))));
assign w54 = (^(6'h11));
assign w55 = {$signed((5'h13)), $unsigned(((27'h1a) !== w76)), $unsigned({(30'h1a), (-9'h1e), w8, (-18'h8), w10, w65, w75, w69, (21'h12), (24'ha), w66, w100, (-6'h1d), w70, w58, (29'h8), (-8'h3), w91}), (-20'h15), (-(w91 ^~ w88)), $signed((w7 ? w100 : (-15'h14))), (10'h16), (^~(-w5)), $signed((^w60)), {(2'h13), w73, (-23'h10), (-27'hb), w74, w1, w83, w69, (-3'h10), (-3'h6), w72, w80, w96}, {w80}, (((-21'h16) ? w90 : (-22'h12)) ? {(-14'h17), (-24'h17), w2, w71, (-17'h1), (9'h16), (31'h6), (8'ha), (-30'h16), w56, (-26'h11), w65, w78, (18'he), (-17'h1d), w68, (-15'h12), w84, (25'hd), w9, (2'h1a), (5'h18), w85, w95, (-20'hb)} : (w75 >= w56)), (9'hf), {(-28'h19), w6, (21'h10), w60, (22'h4), (15'h1d), w80, w100, w65, w85, w64, (-19'h17), (-2'h1e), w9, (17'h7), (10'h15), (9'h6)}, (3'h1d), {(14'h13), (-7'h4), w5, w75, (11'h4), w94, w70, w78}, ((-9'ha) & (~^(-28'hc))), $unsigned((26'h19)), w95, w61, (((16'h17) ? (-19'h3) : (-21'ha)) ? (-17'h1b) : (w58 & w60)), (((26'h5) << w10) ~^ (-23'h3)), w68, ({w69, (11'h17), w80, w99, (-3'h1d), (-6'h5), w4, (7'h11), (-32'h3), w84, w87, w87, (-25'he), w58, w79, (-8'h1b)} ? (~^w66) : (w6 ? (22'h1b) : w65)), w90, ({w82, w65, w85, w3, w66, w5, (25'h7), w59, w84, (2'h17), (10'hc)} ? (+w6) : {(-1'h1c), w63, (-6'h3), (4'hf), w93, w76, (-13'h17), w62, w90, w72, (7'h11), w5, (16'h1d), w93, (11'h8), (-1'h15), (-26'h3), w9, w77, w61, w86, w69, (-3'h7), w5, w80, w93, (-28'h17), (-31'h1a)}), (-29'h12), (-(-24'hf)), ((-19'h1b) || (-21'h12)), (^~$signed(w65))};
assign w56 = {(27'h1b), ((w83 ? (-8'h1a) : w58) * {(-2'h4), (-27'h4), (-24'h3), (-16'h2), (-7'h11), (10'hc), (13'h2), (-9'h8), w93, w72}), ({(-3'h4), w61, (14'h1d), w81, w61, w62, w87, (26'hc), w86, (27'h14), (-5'h1c), w82, (21'h6), (18'h11), (22'h9), (-31'h3), (-19'h16), w1, w73, (-15'h10), w94, w83, w87, (-13'h1), w61, (-29'h0), w72, w85} ? w64 : {(-26'h17), w73, (-25'h3), w70, w95, w68}), ({w78, w10, (-17'h1b), (9'h5), w3, w96, (-1'h1b), (16'h9), (-1'h1d), w62, (20'h8), w73, w80, w80, (-18'hb), w9, w99, (9'h1b), (12'h12), (-24'h1a), w97, (25'ha), (-1'h6), w57, (-9'h1a), w57, (18'h1)} ? w89 : $unsigned(w71)), w70, ((-20'h5) ? {(1'h14), (-12'h1a), w94, w74, (5'h1b), (-7'h10), w87, w68, (-18'h8), (-20'h8), w5, w91, (4'h1d)} : ((2'h4) ? (-24'h1e) : w69)), w85, ({(-15'hc), w95, w92, w69, w65} >> ((7'hf) * w76)), (~|$unsigned(w97)), w90, {(-13'hc), w89, w9, (-11'h1e), (10'h10), (7'he), w84, (19'h1c), (23'h9), (-30'h1a), (23'h16), (20'h1d), (-7'h8), (-6'h3), (15'h14), (23'h18), (-27'h1c), w78, (-18'h2), w94, (31'h1a), w65, w10, (25'h2), w62, w76, w89}, ($signed(w79) ^~ $signed((8'ha))), ((+(-7'h8)) ? (w96 ? (18'hb) : w88) : $unsigned((10'h15))), ({(22'h8), (-2'h11), w61, (22'h11), w70, (12'ha), (-5'h12)} ? (~^(29'h11)) : (^~(23'h10))), (-13'h1d)};
assign w57 = (-8'h8);
assign w58 = ((~&$signed(((w63 == (10'h10)) ? $unsigned(w78) : {(39'h7), w73, (8'h10), w91, w66, (-9'h4), w5, w79, (3'h6), w77, w2, (-29'h1a), (17'h6), w2, (-11'h1d), w86, (-29'h1b), (17'he), (-14'h16), (-5'h15), (-2'h4), w65, (26'h6), w98, (-9'h15), (-8'h1), w87, w66, (17'h6), w100}))) & {((2'h1) ? w66 : (-22'h15)), w2, ((9'h18) ^~ (-25'h8)), (-8'h1c), w67, (29'h3), (w94 ? w60 : (-25'h1)), $unsigned((30'h10)), $signed((21'h6)), (23'he), (w87 >>> w88), (9'h7), $unsigned(w80), w59, (-4'h19), {w80, w88, (6'ha), w79, w10, (5'h2), (-4'h2), (-5'he), (7'hd), w72, (6'h1a)}, (24'h17), w3, ((15'h6) ? w62 : (-22'he))});
assign w59 = ($signed({w100, w82, (20'hc), (9'h7), (-28'hf), (-26'h1d), w87, w88, (21'h1e), (7'h1c), (-10'h0), (31'hb), w70, (-9'h1d), (6'h10), (-24'h3), (-32'h14), (-6'h12), w100, w9, (-25'hf), (22'h1b), (-23'hc), w61, w64, w65, (20'h15), (5'h5)}) < $signed($unsigned({(-25'h1d), (-3'h12), (-1'hf), w79, (30'he), w77})));
assign w60 = (29'h4);
assign w61 = (+(10'h6));
assign w62 = w67;
assign w63 = ($unsigned((w6 >>> (+(w76 ? w80 : w3)))) | (-24'hf));
assign w64 = ($unsigned(w68) ? (9'h13) : {(-9'hb), (+w75), (^~w69), {w87, (-14'h4), (8'h18), w76, w86, w66, w3, w97, w82, w7, w100, (9'hb), (16'h7), w93, (18'h16), (29'h14), w3, (6'h16), (-26'h1), (15'h2), (20'hb), (-12'h1b), w84}, w83, (w66 ~^ w85), ((-1'h6) | w69), (w72 + (-16'h1e)), (-12'h18), (~|w65)});
assign w65 = ((26'h15) + (-13'h2));
assign w66 = ($unsigned(w88) <= (21'h8));
assign w67 = (($signed((3'h7)) ? w1 : ({(-16'h15), (-6'h2), w93, (4'h8)} && $signed($signed((10'h19))))) >> (w77 ? {w3, w3, (-11'h2), w4, (19'hc), w86, (-17'h12), (-28'h12), w98, w68, (13'h18), w77, w3, (-18'h1), w89, (-11'h16), (-20'ha)} : ((w89 < w70) * (w89 | ((-25'h1a) ? (-25'h14) : w5)))));
assign w68 = (-27'he);
assign w69 = {$signed((~^(31'h6))), (8'h11), ($unsigned(w74) ? ((5'h8) ? (29'h4) : w78) : (32'hf)), $unsigned((w71 << (-8'h1b))), w3, ((-7'hb) + $unsigned(w89)), $signed((23'ha)), (31'h1c), (-(w92 ? (-25'h15) : w80)), ($unsigned((-25'h8)) >>> w7), (+$unsigned((-27'h1d))), w2, ((17'h3) ^ {w2, (14'h19), (-30'h2), w81, (18'h16), (19'h2), w86, (1'h1b), (-22'h15), w91, (16'h2), w3, w74, (-3'hf), w9, w76, w7, w5}), (w1 ? w3 : $signed((6'hf))), w1, {(-14'h12), w76, w84, w6, w7, w70, (18'h1d), (-11'he), (-1'h0), w83, (-14'h11), w76, (-8'h0), w93, (30'h13), w1, (-21'hc), w9}, (((7'ha) ? (-30'h12) : (-28'h5)) ? $signed(w98) : (w97 && w74)), ((w76 | w91) ? $unsigned(w93) : $unsigned((-5'h12))), $unsigned((20'h8)), ($signed(w89) < $unsigned((-12'h0))), {w95, (-11'h1e), w83, (-28'h1b), (-15'h8), w92, w95, (-10'h11), w76, w5, w1, (16'h2), w89, w3, (-3'h4), w95, (8'h7), w78, w88, (27'h16), (-30'h19), w89}, (-6'h18), {(-31'h15), (-6'h3), (25'h10), w73, w1, (21'h16), (5'h11), (-24'h5), w95, w96, (-24'h9), (-5'h4), w73}, ((w82 || w87) && (!(10'hd))), w86, {w4, w77, (28'h14), (-8'hd), w8, w87, w79, w6, w74, w79, (-22'ha), w93, (8'h13), w8, w100, (-24'ha), (18'he), w77, w7, w7, w92, (32'h1), w3, (-7'h3), (-9'h12)}};
assign w70 = (-5'h13);
assign w71 = ((w93 ? ((-3'h2) ? ((-22'h1c) << (-5'h2)) : w89) : ($unsigned(w88) ? (~|w74) : {(-28'h1c), w3, w77, w78, (23'h16), (-11'hc), w89, w79, w72})) ^ ((^~$unsigned({w97, (-7'h4), (27'h8), (-9'h1a), w87, (6'h2), w92, w89, w10, w4})) ? $unsigned(w94) : w9));
assign w72 = (-30'hf);
assign w73 = ((12'h1b) < ((~&(+w91)) ? {(-23'h7), (8'h1a), w96, (-25'h9), (-5'h7)} : (-$signed($unsigned(w87)))));
assign w74 = $unsigned((-w78));
assign w75 = $unsigned($unsigned(((-16'h1d) ? (23'hf) : $signed(((-26'h16) ? (9'hc) : (-6'h18))))));
assign w76 = (|$unsigned((((&(8'h1b)) === $unsigned(w1)) != (-4'hf))));
assign w77 = w99;
assign w78 = ({(~|(-22'h4)), (w88 - (13'h1d)), (~&w95), (w3 ? (21'h11) : w99), (+w5), {w93}, w91, (-w8), (|(27'h1b)), (21'h1c), {(10'h1c), (-28'h1c), (34'h2), (7'h1b), (12'he), w6, (10'h1a), w98, (22'h10), (28'h1a), (-16'h1d), w93, (-1'h1e), (-22'hb), (23'h14), w88, w98, (-4'h4), w4, w5}, w86, w81, $unsigned((-14'hb)), ((-26'h12) >> w82), w89, {(-26'he), (-12'h12), w84, (9'h8), w96, w80, (-10'h17), (-23'h0), (-11'h6), w5, w91, w93, w85, (-5'h0), w92, w88, w6, (30'h11), w96, w93, (36'hd), w85, (28'h8), (28'h13), (-18'h3)}, {(28'he), (14'h19), w96}, ((-28'h17) ~^ w85), ((-16'h1a) < (-29'h1d)), {w97, w100, (6'h10), (30'h1d), w5, w97, w89, (7'h7), w81, (22'h2), w96, (20'h19), w99, w3, (-28'h1a), w95, w81, (-6'he)}, (w4 ? (-6'h1b) : (-22'h5)), ((22'h14) ? (-13'h1b) : w94), (w90 ? w93 : w99), (~&w3), {w10, (2'h1e), (16'h19), (25'h7), (-25'he), w85, w81, (-30'h9), w8, (-26'h9), w94, w80, (-10'h2), (10'h10), (-13'h1c), (12'h1b), w83, (31'h4), w5}, w9, $unsigned((-15'h7)), (29'h16)} ? (((w94 >>> w85) ? ((10'h11) ? (31'ha) : (12'h1a)) : w5) & ({(17'he), (9'h18), w93, w4, w90, (-6'h13), (-26'h16), w2, w5, (-10'h4), w5, (-13'hb), (3'hb), w5, (8'h17), w93, w3, (28'h1), w7, (-3'hc), w83, (1'h6), w84, (-21'h8), w82, w82, (3'h4)} << (10'h2))) : w94);
assign w79 = {((~^(10'h12)) != (w2 >= (12'hf))), {w4, (-9'h5), (18'h16), (18'h7), (24'h11), w83, w82, w3, (3'hc), (2'h19), w82}, ({(27'h1e), w95, (25'h1c), (-26'h17), (14'ha), (-23'h16), (7'h7), w95, (-14'h4), w81, (-19'h4), w90, (-13'hf), (2'h19), w2, w99, w88} & {(-29'h13), (-7'he), w84, w5, (-22'h11), (10'ha), (-11'h1e), w92, (-30'h19), (-1'h11), w9, (-20'h4)}), (~|(&(3'h12))), w84, (^((16'h12) <<< (-28'h1a))), w85, (((6'h17) ? (16'h17) : w94) ? (w5 & (15'h1a)) : (w86 != w85)), w8, w89, w89, w88, ((w80 ? w7 : (28'h17)) ? (^(7'h10)) : (!(26'hf))), ($unsigned((11'hf)) ? {w83, w4, w96, (-12'h1), (-29'h1e), w10, (-17'h6), (-11'h2), (-5'h0), (3'h1c), (15'h3), (2'ha), w5, (8'h3), w82, w96, (-32'h2), w80} : (~&w4)), $unsigned((w10 ~^ (13'h15))), (30'h10), (~^(-15'h13)), {w98, w4, w99, w8, (5'h18), w84, w7, (-20'he), w85, (26'h7), w100, w93, (-16'h1a), w6, (27'h3), (-15'h8), w82, (28'ha), (18'h8), w2, (-1'he)}, (((-15'h9) ? w6 : w97) | w93), $unsigned((w87 ~^ w4)), $unsigned({(-25'h5), w92, (-4'h1e), w9, w10, (17'h1c), (1'ha), w2, w98, (-9'he), (29'h3), (-2'h6), w92, (-20'h8), (5'h1c), w100, w94, w5, (-15'h16)}), ({w3, (-19'h1a), (-22'h5), (-4'h9), (-17'h19), w80, w4, w85, (-13'h1c), (12'h15), (-22'h1), (2'hb), w85, w7, (-3'h4), (32'h1c), (-26'h4), (-16'h1d), w97, (25'ha), (18'h7), (23'h8), (3'h15), (10'h13), w99, w9} !== w8), (26'hd), (|((28'h13) * (20'h8))), {w10, w98, w80, w10, w10, (-1'h1d), (16'h1d), w91, (1'h8)}, {(4'ha), (23'h1e), (23'h3), (16'h1a), w83, (-28'he), w6, w90, (5'h5), (-4'h1e), w83, (-31'h6), w96, (-22'hc), (-22'h5), (-25'h2), (-32'h0), (-22'h14), (-14'h1a), (26'h12), w3, w88, (8'h6), (22'h3), w84}, {(-5'h15), (26'h1a), w1, (5'h6), w95, (18'he), w87, w85}, (((16'h1d) < (16'h3)) | (~|w3)), ({(23'h2), (16'h3), (19'hc), w9, (-19'h14), (-18'h1b), w99, (-22'h15), (-22'h1a), (-15'hf), w100, (26'h1e), (-17'h18), w8, (23'hb), w90, w96} ? (!w85) : (~|(-24'h4)))};
assign w80 = (-23'h1b);
assign w81 = (-23'h5);
assign w82 = $unsigned({w100, (w10 <= w9)});
assign w83 = $signed(((((4'h19) >> (16'h1a)) ? (5'h10) : (|w87)) ? w6 : w98));
assign w84 = w4;
assign w85 = ((7'hb) >>> ({(-16'h13), w1, (23'h6), w95, w9, w10, (-3'h18), (-7'h18), (-18'h1d), (18'h6)} ? (^~w4) : (|((w90 | w93) == (24'h3)))));
assign w86 = (w8 ? {(w92 * w90), {(-18'h12), (-14'h0), w6, w3, (17'h6), (1'h1), (-19'h15), (-18'h12), (-17'hb), w92, (-26'h1a), (16'h11), w94, w96, w90, (24'h5), w95, w97, (-19'h17), w100, (-28'h1d), (25'h9)}, {(-21'h4), w6, (16'h12), w91, w97, w94, w95, (-9'h8), w1, (-1'hc), w7}, w93, (15'h12), (8'h10), w3} : (-2'h11));
assign w87 = (&(((w4 ? w90 : w4) ? (w95 ? (-17'h10) : w93) : (+(18'h8))) ? w91 : ((((-14'h3) > (20'ha)) | $unsigned((-18'h0))) <= w90)));
assign w88 = (((-15'ha) ? ($signed({w99, (20'h16), (-25'h1)}) >> (((-26'h15) ? w3 : (-23'h16)) <= (-18'h7))) : (-6'h1b)) * ({(15'h4)} ? (~^{w10, (-13'h1b), (-1'h19), (-10'h7), w100, w7, w5, (-4'h1a), (27'h13), w94, w9, w97, (15'h1a), (-15'h2), w7, (29'h9), w5, (19'h10), (28'h5), w90, w100, w96, (26'h3), (10'h19), (2'h12), (26'h12), w91, w3}) : (^~(w3 !== $unsigned((-5'h1e))))));
assign w89 = w2;
assign w90 = (~&(+{w93, (29'h19)}));
assign w91 = (($unsigned((27'h10)) ? (-16'h1e) : {(17'h3), (-11'h12), w93, w96, (-1'h1b), (-23'h8), (-21'h18), (-27'h8), (23'h13), w9, w98, w94, (-24'h4), w5, w92, w9}) ? ($unsigned((w97 ? (1'h19) : w7)) ? ($unsigned((30'h14)) ? (|(30'h7)) : (w96 ? w93 : w5)) : $unsigned((-9'h10))) : {(w96 & w98), $unsigned((8'h14)), {w2, (6'h16), (-16'hd), w4, w3, w10, (-11'h7), w5, w10, (-21'h1d), (-23'hb)}, (w10 ? (14'h14) : (27'h16)), $unsigned(w7), {w5, w93, w2, (5'h7), w6, (6'h5), (-3'h5), (26'h2), w93, w96, (1'he), (-20'h3), (-2'h1a), w9, (-16'h1b), (5'h17), w5, w3, w8, w95, (-23'h5), w3, w92, w97, (-29'h1c), (-7'h10), w92, w95, w1, w5}});
assign w92 = $unsigned((-22'h2));
assign w93 = {($signed(w3) <= w8), ({(-24'h7), w10, (-26'h6), (-18'h15), (24'he), (26'ha), (27'hd), (13'h19), (25'h10), w8, (-10'h1a), w100, (-3'h3), w96, (-28'h3), w9, w98, w98, w8, w100, (-17'h1d)} >> (|w100)), $signed({(28'he), (-28'h15), (22'h6), (-30'h18), (18'hb), w97, w3, (-18'h13), w5, w7, w3, w98, w100, w95, (-15'hb), w5, w96, w7, w7, (-4'h14)}), (~^$unsigned(w100)), (-3'ha), ((22'hb) & w2), ((w3 ? w5 : (-3'h8)) ? w100 : (~&(-16'h12))), (-18'h4), w98, ((w4 && (-20'h7)) | $unsigned((28'h1a)))};
assign w94 = ((-10'h16) ^ w98);
assign w95 = ((1'hf) == ((~^$signed((w7 << (-9'h16)))) ? $unsigned(((-19'h14) ? w8 : (28'h11))) : (|{(26'hc), (18'ha), (27'hd), (16'hd), w96, w10, (24'h2), w98, w96})));
assign w96 = (((~|((w8 ? w1 : (26'hf)) ? (17'h16) : ((22'h7) | (-12'h2)))) || {w6, w99, (-20'h5), w8, (-14'hf), w98, (26'h6), w9, w99, w99, w8, w99, w9, w10, (-17'h19), (-24'h6), (-25'h3), w3, (-26'h1d), (22'h16), (-18'h19)}) == {(-5'h4), {(-16'hf), (11'h2), w1, w9, (14'h15), w1, (5'h5), w100, w6, (15'h8), w8, (9'h1d), (31'h4), (-26'h19), w97, (-23'h1e), (-27'h1c), w98, (-14'h19), (-22'h17), w9, w3, (18'h6), w97, w7, w98, w5, w7}, $unsigned(w99), (w8 <= w2), ((17'h7) ? (-5'hd) : (30'h1a)), (&w5), (1'hd), (w1 == (10'hb)), (w4 ? (14'h10) : w1), (w100 ~^ (14'h2)), ((20'h2) ? w2 : w100), ((-7'h15) ^~ (25'h1e)), (w4 ^~ (-21'h13))});
assign w97 = (~^({w5, w7, (-17'h18), (30'hf), w1, (-3'h14), w6, w98, (-10'h12), w2, w100, (10'h3), (21'h9), w4, w6, w5, w99, w7, w1, w100} ? {(-14'h7), (-28'h16), (25'h1b), (14'h7), (26'h1d), (9'h14), (-22'hc), (6'h1d), w10, (5'h8), w10, (5'h1b)} : $unsigned($signed(((-29'h12) <= (-19'h14))))));
assign w98 = w99;
assign w99 = ($signed((29'hd)) > $unsigned($signed(((1'h13) >> (w100 ? w5 : (-9'h9))))));
assign w100 = w7;
assign y = {w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100};
endmodule
