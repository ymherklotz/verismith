module test_module(y, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10);
output wire [1472:0] y;
input wire [23:0] w1;
input wire [20:0] w2;
input wire [1:0] w3;
input wire [29:0] w4;
input wire [23:0] w5;
input wire [22:0] w6;
input wire [20:0] w7;
input wire [26:0] w8;
input wire [3:0] w9;
input wire [8:0] w10;
wire [10:0] w11;
wire [27:0] w12;
wire [2:0] w13;
wire [24:0] w14;
wire [1:0] w15;
wire [6:0] w16;
wire [2:0] w17;
wire [21:0] w18;
wire [9:0] w19;
wire [27:0] w20;
wire [8:0] w21;
wire [9:0] w22;
wire w23;
wire [23:0] w24;
wire [2:0] w25;
wire [13:0] w26;
wire [28:0] w27;
wire [18:0] w28;
wire [29:0] w29;
wire [28:0] w30;
wire [12:0] w31;
wire w32;
wire [21:0] w33;
wire [9:0] w34;
wire [20:0] w35;
wire w36;
wire [27:0] w37;
wire [22:0] w38;
wire [26:0] w39;
wire w40;
wire [5:0] w41;
wire [21:0] w42;
wire [10:0] w43;
wire [14:0] w44;
wire [26:0] w45;
wire [16:0] w46;
wire [23:0] w47;
wire [26:0] w48;
wire [2:0] w49;
wire [24:0] w50;
wire [8:0] w51;
wire [8:0] w52;
wire [27:0] w53;
wire [4:0] w54;
wire [12:0] w55;
wire [26:0] w56;
wire [18:0] w57;
wire [18:0] w58;
wire [27:0] w59;
wire [14:0] w60;
wire [6:0] w61;
wire [21:0] w62;
wire [28:0] w63;
wire [17:0] w64;
wire [4:0] w65;
wire [19:0] w66;
wire [28:0] w67;
wire [7:0] w68;
wire [21:0] w69;
wire [16:0] w70;
wire [14:0] w71;
wire [10:0] w72;
wire [7:0] w73;
wire [9:0] w74;
wire [26:0] w75;
wire [15:0] w76;
wire [22:0] w77;
wire [21:0] w78;
wire [16:0] w79;
wire [7:0] w80;
wire [19:0] w81;
wire [28:0] w82;
wire [6:0] w83;
wire w84;
wire [13:0] w85;
wire [13:0] w86;
wire [21:0] w87;
wire [25:0] w88;
wire [26:0] w89;
wire [24:0] w90;
wire w91;
wire [26:0] w92;
wire [3:0] w93;
wire [16:0] w94;
wire [18:0] w95;
wire [23:0] w96;
wire [11:0] w97;
wire [10:0] w98;
wire [26:0] w99;
wire [9:0] w100;
assign w11 = (~|$unsigned((w49 > $unsigned((w31 < (17'h7))))));
assign w12 = ({w65, (w41 == w52), ((7'h4) ? w44 : w3), ((7'hf) ? w59 : w69), $unsigned((19'h1)), {w95, (20'hb), (24'h3), w92, w44, w45, w25, (-27'h11), w58, w76, (16'h10), w35, (-29'ha), (-16'h18), w97, w28, (-7'h2), (-18'h6), w69, (4'h8), (-5'h15), w63, (26'hf)}, w27, (-19'h1d), (^w50), {(-7'h2), w53, (-28'hb), (-3'h1b), (-23'h6), w66, (-26'hf), w82, (-4'h11), (-2'hc), (-6'hc), w37, (27'he), (20'h3), w50, (-21'h18), (30'h3), w25, w54, w53, w55, w40, w34, (28'h7)}, {(-14'h1c), w77, (-25'h16), w56, (-27'h1), w40, (27'h19), (-24'h1), w33, w46, w41, w70, w62, w89, w9, w71, w31, w30, (-1'h16), (-10'h1e), (-3'h0), (-25'h16)}, {w91, w79, (-27'he), w9, w73, (-6'h10), w5, w76, w55, (7'h16), w38, (-12'h11), w53, (12'h18), (-25'h4), (-28'h1e), w54, (14'hf), (-15'h7), w98}, ((31'h19) ? (-33'ha) : (8'h1)), (w96 ? w52 : w49), {(-15'h11), (-26'h2), (21'h18), w87, w63, (-28'h1), (-30'h1), w54, (-22'h1e), w90, (-31'h0), w9, w87, w84, w22}, $unsigned((-32'h3)), (!(-10'h1))} !== {$unsigned((-3'h13)), ((-4'h16) & w78), w56, {(28'h3), w26, w87}, ((11'hb) != (-24'h14)), (|(-31'hc)), (-5'hf), $unsigned((-27'h1c)), $signed((19'h4)), w42, (+(-24'hf)), w4, $unsigned(w6), (|w83), $unsigned((-11'hc)), w1, (-(-10'h0)), $unsigned(w20), w74});
assign w13 = {{(-6'h2), w70, (-13'h17), w5, w4, (17'hb), w7}, ({(-6'h1c), w61, w47, (2'h10), w2, (4'h8), w31, (12'h14), w65, w61, (-26'h18), w34} ^ (w47 <= w26)), w62, $unsigned(((17'h1e) == w76)), (6'h11), (-30'h14), (20'h19), $unsigned($unsigned((33'h17))), $unsigned(w50), w76, {w78, w48, (-22'hb), (18'h6), (-30'h1), w92, w97, (8'h6), w89, w62, (-23'h9), (11'h2), w20, w81, w54, (12'h10), (16'h4)}, {(-28'hf), (27'h13), w4, w44, (25'h12), (-15'h12), (7'h3), w100, (-17'h11), (7'h1a), w64, (-9'h10), w24, w51, w63, w81, (12'h8), (-4'h1b), (-14'h3)}, w36, ((w70 | (-23'h17)) ^ (!(26'he))), (11'h15), (-30'he), {(-10'h1)}, (|w51), (~^w5), (5'h1b), ($unsigned(w45) ~^ w78), (((-27'h14) >> (-30'h3)) ? $signed((-19'he)) : ((25'h9) | (14'hd))), w54};
assign w14 = ((^($unsigned((30'h1d)) ^~ (^~w68))) !== w42);
assign w15 = (-13'h8);
assign w16 = ({(-5'h16), (20'hd), $signed((22'h10)), w28, w45, {w23, (-20'h13), w67, (30'h12), (-14'he), w71, (-24'he), (-28'h16), w7, w50, (-12'h15), w58, (25'h13), (8'h4), w100, w79, w19, w73, (-30'h4), w54, (20'h4), w24, w82, w97, w74, (-12'h1), (18'hd), (-28'hb)}, (w79 ? (6'h16) : (16'h10))} || (^(17'he)));
assign w17 = ($signed((~&((~&(28'h5)) << ((-4'h19) ? w59 : w51)))) ? $signed({w94, (9'ha), w65, (17'hd), (-9'h11), (-22'hb), (-22'h8), (-21'h11), (9'h16), w36, (13'h5), w9, (-18'h18), w35, w29, (-11'he), (-31'h1c), w62, w75, (-2'h19), (27'h9), (-28'h7), (28'h1d), w23, w67, (12'h11)}) : (26'h6));
assign w18 = w47;
assign w19 = w61;
assign w20 = ((-10'h1d) & (~&{(-13'h2), (-2'hb), (-9'h1d), (5'h4), w50, (16'h3), (-14'h19), w32, w98, w36, w22, (19'h5), (-10'h19), w79, w22, (6'h6), (-1'hb), (-3'h8), (29'h6), w59, (-23'h9), (-27'h10), w29}));
assign w21 = w49;
assign w22 = w64;
assign w23 = (21'h1c);
assign w24 = ((({(-19'hb), w81, (12'hf), (25'h18), (10'h7), (27'h3), w56, w31, w2, (-30'h2), w37, (28'h15), (20'h12)} ? w84 : {w41, w36, w98, w50, (22'h8), w81, w49, w96, w98, w50, w64, w62, (20'hf), w40, (27'h9), (20'ha), w84, w42, w10, (29'hd), w40, w1, (25'h8), w7, w90, (18'h2), w68, (28'hd)}) ? w87 : ($unsigned(w51) <<< $signed((16'h2)))) ? {{(-2'h0), w59, w45, w52, (27'ha), (-22'h1c), w78, (21'h6), w89, (24'ha), w87, (-30'h8), w8, w8, w25, w32, (-20'h2), (3'h11), w86, (-17'h1a), w73, w100, w100, w77, w71, w64, (-15'he)}, $unsigned(w32), {(30'h1), w95, w86, w52, w59, (24'he), (-27'h1b), w69, w37, w75, (15'h11), w60, (-21'h5), (-11'he), w40}, (-w95), (-26'h2), (-4'h11), w5, ((10'h13) && w60)} : $unsigned((~^(((14'h8) ? w50 : (16'h18)) >>> {(-11'h1a), (12'h8), w70, w49, w50, w3, w74, (-13'h4), w41, (-31'h1d), (29'h7), (-22'hc), w90, (14'he), w86, (28'hd), (21'h6), w81}))));
assign w25 = (^~{(15'hf), (w85 ? w59 : (-7'hb)), (~^(-12'h17)), (-29'h0)});
assign w26 = $unsigned({w57, ((-17'h18) < w93)});
assign w27 = w59;
assign w28 = (-4'h15);
assign w29 = ($signed(w93) >= (-(w62 ? w4 : {w69, w8, w100, (-8'h12), w66, w42, w100, (-8'h10), w69})));
assign w30 = {((-1'h1b) ? w61 : (10'h6)), ($unsigned(w86) ? ((1'h1e) < w75) : w66), ({w69, (-21'h4), (-7'h7), w39, (13'h11), (-9'h13), w55, w46, w93, (6'h7), (22'h1b), w58, w54, (15'h1b), w83, w1, (6'h15), w51, (-5'h10), (12'h12), w40, (-3'h8)} ? {(12'h10), (4'h4), w61} : (-30'h5)), {w93}, w69, ({w84, (-12'h1e), (22'h8), w65, w53} ^ (^w100)), $signed((w9 ? (-29'h1c) : w31)), $unsigned((w59 ? (-6'h2) : w93)), {w52, (10'h16), w41, (-17'h16), w51, w98, w1, w54, (16'he), w82}, (!(3'h14)), $unsigned($unsigned(w68)), w66, (-29'h5), $unsigned((w4 ? (-15'h9) : w45)), (11'h3), ((16'hd) < (-8'h2)), w68, (23'h1e)};
assign w31 = w37;
assign w32 = (^~((-1'he) ? w75 : {w73, w71, (-1'h14), w62, (-36'h1b), w57, (-5'h6), (-3'h1d), (24'h19), (-12'h14), (-17'h15), (4'h19), (-26'he)}));
assign w33 = $signed((w68 | (-13'ha)));
assign w34 = $unsigned($unsigned((14'h1d)));
assign w35 = (|($signed((23'h16)) ? $signed(w39) : ((6'h8) ? (w54 ? w73 : w69) : (&(-15'h10)))));
assign w36 = $unsigned(($unsigned((w70 > (~&w74))) ? w47 : {(19'h10), w1, (5'hb), (20'h1c), (15'h1), w46, (-25'hf), (-6'h18), (-27'h13), w94, (3'h18), w54, w75, (24'h1b), (-11'h14), (14'h7), w82, (-11'hb), w98, (-19'ha)}));
assign w37 = (+(|((-27'h5) * (-32'h13))));
assign w38 = $unsigned(({w71, (-9'h8), w42, w62, (13'h9), (29'h8), (-24'h1c), w57, w8, w73, (-13'h2), (-1'h2), (2'h16), (9'h16), w79, (-10'h7), (10'ha), (-15'h19), (27'h16), w82, w52, w84, (-19'h14), w10} ? ((^(3'h6)) ? (-19'ha) : w91) : $unsigned(w53)));
assign w39 = {(w3 == w57), w62, (17'h15), (-(w8 ? w67 : w57)), (w51 - $unsigned((-29'h13))), w67, $unsigned((&w99)), (^(~&w9)), (((23'h1b) === w55) ? ((28'ha) ? (19'h16) : (3'h8)) : (+w86)), {w60, (13'h5), (-15'he), w7, (12'hb), (-8'h0), (14'h4), w79, w74, w56, w62, w7, w1, (-19'h11), w2, (31'h16), w95, (14'h5), w67, w53}, (~^$signed(w80)), (~&w89), (10'h17), (12'h7)};
assign w40 = $signed({((5'hd) !== (2'hd)), $signed((-30'h1d)), (w52 <<< w84), ((15'h10) ^ (-31'h9)), {(1'hb), w85, (-17'h15), w58, w87, (7'h6), w50, w85, (-2'h2), (28'h8), (22'hf), (34'h17), (22'h15), w70, (22'h3), (15'h1e), (-25'h3), (-9'h8), (-2'h1a), w42, (-1'h2), w95}, ((-18'h1a) < (30'h7)), {(-8'h7), (-16'h1b), w79, w50, (-4'h1), w53, (-7'h11), (20'h16), w91, (18'h6)}, {w83, (-25'h1e), w2, (11'hb), w61, w90, (-6'h1)}, $unsigned(w81), (w92 <= w86), (!(-26'h11)), $unsigned(w89), (w73 ? (-7'h13) : (-16'h19)), ((-14'h13) ? w55 : w63), {w97, (-22'h19), (3'ha), w47, (-1'h19), w98, (19'hb), w68, (-13'hb), w61, (5'h10), w1, w57, w63, w74, (-30'h13), w50, (-16'h1e), (-8'hf), (-21'h1c), w46, (-9'hb), w86, (-22'h6), w84, w90, w96, w84, (-24'h1)}, (~&w74), w89, (|(19'h19)), ((-16'hf) != (-10'h8)), (w86 && w74), (w55 >= (13'h1c)), (w46 < (-30'h14)), {w50, w67, w92, w54, w65, (-18'h9), (29'h2), (-17'h1b), (-11'h0), (-18'hd), w86, w4, (14'h8), (-28'h18), w88, w5, w51, (-30'h12), (-18'h12), w41}});
assign w41 = $unsigned(((-24'h1e) == (!w79)));
assign w42 = (!{(11'h1e), (w53 ^~ (-18'h7)), {(-22'h5), w59, (5'h17), w64, w81, w65, w98, (2'h12), w6, (29'h1), (2'h14), w47, (19'h17), (-13'h13), w54, w79, w2, (-4'h8), (-14'h1a), w92, (6'h1b)}, w59, (w65 >> w98), $unsigned(w94), $signed((14'h1b)), w10, ((27'h6) >> (-32'h19)), (w67 >> (13'hf)), {(19'h18), w1, w70, w71, w83, (20'h1a), w85, w2, (6'hd), (21'h1d), (15'h16), (-11'h18), w80, (-13'hb)}});
assign w43 = $signed({$signed(w1), (-w51), (-(-10'h13)), (&w60), $signed(w78), $signed(w8), (9'h3), w7, {(-11'h4)}, ((8'h16) != (-30'h3)), ((-6'h16) ? (-1'h0) : w50), ((1'h19) <= w83), $unsigned((-9'h18)), (!(3'h7)), (w45 ? (-32'h0) : w62), w67});
assign w44 = (+($signed(((17'hd) >> w5)) != (^~(25'h18))));
assign w45 = w89;
assign w46 = $signed({(-15'h2), {w93, (-24'h0), (-17'hd)}, {(26'h1d), w55, (-23'h0), (1'h4), (15'hd), (-15'h1e), w54, (11'h2), w6, (-20'hf), (2'h16), w100, (20'h1a), (7'h5), (5'h17), (-2'h13), w97, w56, (-6'h4)}, $unsigned((31'h1)), ((-31'hb) > (-33'ha)), $unsigned((-8'h11)), (^w95), (-w4), (29'he), $signed(w48), (|w68), (18'hc), {(-29'h10), w2, w9, (15'h1b), w77, (-28'ha), (17'h15), (-24'he), (-28'h0), (-30'hd), w47, (-36'h5), (-29'h1e), w81, (-1'h1d), (-1'h8), (32'h8), (17'h9), (4'h9), (-32'hf), w9, (19'h10)}, w78, (~^(-20'h17)), ((21'h12) ? w86 : w5), (w1 >= (1'h1c)), w68, $signed((22'h19)), (w5 <<< (-13'h11)), w63, {w75, (-12'h1c), (-11'h0), (-30'h1b), w8, w70, (-5'h8), (-27'h0), w91, w65, (15'h16), (7'h19), w77, (-32'h18), w2, w94}, (|w57), ((13'h1d) != (-19'h13)), (-3'h17), w5, w76, $signed(w57)});
assign w47 = w7;
assign w48 = ($signed({(-3'hd), (16'h13), (33'h1c), w69, (29'hb)}) ^ {{w58}, (10'hb), (-15'h1b), w5, (~^w73), {w75, (14'h18), (13'h18), (-25'hc), w5, (-32'h1b), (5'hb), w66, (1'h1b), (6'h7), w60, (-20'h13), (20'h1d), (-19'h17), (-12'hd), (18'h1c), (26'h12), w97, (-14'h0), (24'h10), (-6'h9), (-10'hd), (26'h15), w79, (-10'h10), w77, (10'h2)}, ((-14'h1) ? w63 : w87), w59, {w73, (-30'h16), w49, (-12'h1e), (22'h12), w50, (-16'hb), (-4'h8), w75, (8'h17), w97, w93, (-19'h13), w6, (4'hb), (-18'h1d), (-5'h17), (-8'h0), w71, (-3'h1), w64, (-28'h17), w80, w97, (9'he), w68, w71, (-28'hc)}, $signed((-17'h6)), $unsigned(w97), (w93 ? w1 : w70), $unsigned(w72), w77, {w84, (-23'ha), (24'h1b), w87, (-29'h8), (-8'h4), w10, w59, w76, (-20'h14), w96, (-10'h9), w2}, $unsigned(w86), (-9'h1d), ((3'h15) ? w94 : w53), (w90 - (-16'h15)), $unsigned((27'h7)), $unsigned((-4'h16)), $unsigned(w9), ((-27'h1b) ^ w98), (w9 >= w77), (+(29'h8)), ((-18'h1b) <<< w98), ((-12'h19) < w52)});
assign w49 = {$signed((~^w4)), (-17'h1), {w73, w85, (14'h1), w62, (-15'h16), w73, w80, w95, (-31'h14), w57, (-4'h1c), w73, w77, w64, w79, w76, (17'h13)}, w73, w94, (!$signed(w83))};
assign w50 = w73;
assign w51 = (&w73);
assign w52 = (|w82);
assign w53 = (({w78, (14'h1c), w95, (-7'h18), (26'hd), w5, (32'h12), (9'h1d), (-10'h12), w65, (-22'h17), (-27'h17), (32'h11), (-8'h0), (8'h4), (-8'ha), (-11'hd), w97, (25'h6), (12'h3), w90, w76, w9} ? $unsigned(((-7'h15) ? (-21'h1a) : w91)) : w60) >> ((|(~^w74)) ? {(-9'h0), (26'h7), (26'h18), (17'h7), (-22'h5), (-18'h3)} : (w68 == (w4 ? w9 : (32'h18)))));
assign w54 = (~^((({(-27'h13), w63, w6, (-4'hd), (20'h1e), (-20'hd), (-22'h16), (27'h7), (14'h13), (-21'hc), w74, w100, (-5'h19), (-16'ha), (-31'h14), w96} <= (34'h19)) ? (&{w74, (29'h1b), (-17'h1a)}) : (w74 <<< (!(10'h1b)))) || w60));
assign w55 = ({(-w85), $signed((17'h19)), {w4, (-19'h10), w63, w84, w79, (-24'h14), w67}} ? (2'h10) : {{(-25'h13), w79, w67, w3, w83, w85, w62, (30'h18), (-27'h1a), w1, w64, w60}, w83, (~&(21'h12)), (-14'h1b), {w76, w57, (-22'h1), w72}, ((26'h8) ^ (30'h13)), (w90 ? w65 : w89), (~^(20'h8)), ((3'h19) ? (-27'h3) : w63), {w89, (15'h16), w100, w5, w93, (29'h18), (16'h7), (-30'h1b), (-1'h1e), (-18'h10), (-9'h8), w7, (18'h7), (7'h16), w98, w67, w99, (-1'h19), (22'h7), w68}, ((29'h1a) != (-23'h0)), (+(23'h4)), w61, (w84 == (-3'h2)), (w66 != (20'h1d)), (w72 === w84)});
assign w56 = $unsigned({((15'hd) ~^ (23'h4)), {(-10'h17), (24'h11), (9'h3), (12'h9), (7'ha), (20'h1b), w80, w83, w66, w71, (16'he)}, (-w69), ((6'hf) ? (11'hc) : (-2'h5)), $unsigned((13'h14)), ((-27'h13) ? w92 : (26'hb)), (10'he), (12'h16), (-12'hb), (8'h1a), (-29'h1c), (-(5'h2)), (w99 + w59), $unsigned((-8'ha)), (^w70), (17'h19), (+w8), w97, (-8'h1d), (-w88), $signed(w85), {(-9'h10), (30'h1c), (5'h16), w83, (1'h7), (14'h11), (5'h2), (-10'h3), (-21'h17), w83, w64, w99, w80, (3'h11), (22'h17), (-28'h13), w70, (21'h1b), w80}, {(23'h1d), w87, (16'h11)}});
assign w57 = (12'h7);
assign w58 = {((w65 ? (-13'h12) : w66) ? (w79 ? (8'h1) : (-4'h5)) : ((-26'h15) ? (28'h6) : w83)), (27'h1c), (17'h10), (((-22'h13) + w61) ? ((8'h15) ? (-3'h1c) : w90) : w4)};
assign w59 = (~&($signed(((w9 != w85) >> (-19'h12))) & $unsigned($unsigned((-w80)))));
assign w60 = {(29'h15), ((-20'h3) ? (6'h14) : $unsigned((-27'he))), ({w65, (27'h12), w99, w91, (23'h1b), w90, (26'h10), w94, (-14'h1a), (-14'hb), w77, (-8'h1c), w69, w99, (-6'h2)} ? $unsigned(w75) : w71), w98, (-30'hb), {(23'hd), w70, w65, (21'h9), (30'h3), w2, w70, w3, (-22'hb), (-4'h1e), (21'h1b), w68, w79, w90, w65, (1'h1c), (-25'h17), w67, w7, w89, (-22'h4), (18'h12), w67, (-14'hc), w1}, $unsigned((5'h13)), w78, (w7 ? ((17'h17) ? (-27'h4) : (-27'h18)) : w84), (-28'h17), (5'h16), $signed((~&(-18'hd))), ((w95 <= w86) <= {w95, (29'h1c), w93, w93, (-19'h4), (-28'h13), (-7'h16)}), ({(-6'hb), (-7'h15), w75, w91, (-7'hb), (-16'hb), (-9'h6), (-21'h0), w8, w2, (5'h1c), w92, (6'h6), (24'h17), w64, (18'h1d), w65, w4, w77, w65, (24'h1d), w72, (-8'h1b), w8, (2'h16), (2'h6), (-6'h17), (-3'h0), (-15'h1d), w79} ? (!w6) : ((1'h3) ? w97 : (-4'hd))), (-6'h8), (~&w6), w83, (18'h2), w2, (+{(-14'h14), w82, (25'hb), w68, (-20'h19), w5, w10, (17'hd), w72, (-4'h3), (9'h10), (-24'h16), (5'h10), (10'h18), (9'h19), (4'h13), w88, (-16'h17), w4, w2, w9}), (31'h19), w90, (-16'h16), $signed(((-9'h1b) ? w99 : w5))};
assign w61 = ($signed({(-11'h1d), (22'h4), w67, (1'h8), (-15'h10), (24'he), (17'h2), w73, w2}) ? ({(-24'h1e), w84, w88, w85, w80, w71} ? w94 : w62) : ({w81, w5, (23'h2), (-8'h13), (25'h1c), (-19'h1a), (3'hb), (-11'h1e), (8'h4), (-1'h1a), w7, (30'h14), (-10'h12), w80, (12'h17), w74, (5'h16)} ? ({w86, (13'hd), (24'h19), (21'h14), (-33'h1d), (26'hd), w2, (12'h10), (29'h4), w84, (-17'h17), w7, w63, w99, w91, w85, w90, w93, w69, (-30'h3), (3'h6), w94, (20'h7), w79, w73, w83, w97, (-2'ha), (9'h4), w8} ? {(5'h2), (20'h1e), (17'h14), (-9'h7), (24'h8), w64, (-5'h8), (6'h5), (12'h1e), w77, (31'h8), (-7'hc), (-6'h12), (24'h1e), (6'hd), w5, w83, (3'h2), (-12'h8), (-4'ha), (-4'h1e), (28'h10), w3, (-18'h13), (14'h13), (-7'he), w69} : (w87 | w2)) : (-28'h5)));
assign w62 = {(((4'hd) || (-27'hc)) ? ((11'h12) ? (22'h1a) : w6) : (22'h1a)), (^((-16'h2) << w1)), w91, (-20'he), (29'h5), (w73 <<< w3), (7'h1e), {(-11'h12), (8'h1), (11'h13), (20'h12), (29'h7)}, {(-21'h0), (3'h1c), (-10'hd), w87, (-5'h12), (-2'h16), w64, (31'ha)}, w98, (((30'h16) + w76) >> w93), (w97 ^ (w64 <<< w73)), ($signed((-1'hf)) << (w63 != w81)), ((&(12'he)) ? (w3 < w80) : (w77 <<< w72)), ((!(25'hb)) ^~ (^(-10'h12))), ((~|w86) ? w68 : w75), w71, w72, {w67, w72, (-8'h10), (21'h1b)}, (-{w8, w87, w86, w93, (18'h1)}), ((6'h19) - ((-20'h6) ? w65 : (-4'h19))), w83, w75, w77, ({(26'h17), w82, (1'h7), (18'h14), (-10'h5), w91} != $signed((-27'h17))), ((w95 >= w2) & w8), (^(2'ha)), (26'hd)};
assign w63 = (-27'hc);
assign w64 = $unsigned({(16'h8), (^w9), w99, (!w67), (-31'h14), ((22'hc) ? (-27'h13) : (26'h6)), {w91, w67, w98, w90, (3'h12), (11'he), (2'h3), (-30'h9), w68, (15'h5), (4'h14), w3, (19'h16), w6, (-26'hb), (-12'h1a), (28'h17), (26'h14), (29'h9), w66}, (28'h1e), (~|w87)});
assign w65 = {((w83 ? w10 : w68) && w93), ({(21'hc), w6, w89, (17'ha), w71, (23'hf), (16'h14), (-20'h1b)} >= ((-3'ha) ? (-5'h16) : (-5'h1d))), (8'h3), ((~^w10) && w92), $signed((w82 ? w8 : (7'hc))), {w79, (-24'hb), w93, w80, (-15'he), w94, w79, (13'h6), (9'hf), w66, w82, w83, w89, w96, w88, (4'h6), (29'h8), w94, w98, w77, (-33'h6), (-8'h3), w84, (6'h4), (-18'h1d), (-2'h6), (27'h1), w7}, {w85, (-7'h7), (19'hf), w84, (-21'h1c), (-6'h4), (-4'h6), (28'h17), w76, w79, (12'h17), (20'h1b), (24'h2), (9'h14), w71, w9, (24'h15), w1, (-30'hb), w10, (25'h3), (-26'h5), (-14'hb), w2, (30'h16), (-7'hc), (-7'h18)}, w88, ((-33'h5) >= (-1'h12)), $signed(w78), ((19'h12) ? {w87, w100, w98, (19'h8), (11'h4), (-15'h11), (-11'he), w5, w70, w68, (25'h1a), (24'h9), w77, w74, (4'h14), w10, w81, w2} : (w91 ? (26'hb) : w68)), (~&(+(-27'hf))), (31'h2), ((-w93) << (8'h15)), (!(|(30'ha))), $unsigned($unsigned((-22'h2))), w73, ((w74 - (-6'h15)) ^~ {(14'h1d), w93, (-4'h4)}), ((w93 ? (5'h1a) : w89) ? (^w84) : $unsigned(w9)), w81, {(-15'h12), w9, w77, (-23'h11), (-5'h1a), (-22'h1b), (-2'hc), w74}, ((|w89) ? {(-1'h0), (-31'hf), w83, w96, (-20'h14), (10'h1e), (8'hd), (-4'h3), (13'h18), (-20'h2), (-11'hb), w87, (-1'h5), w95, w88, w5, w4, w70, (12'h1a), w79, w91, w99, (-27'h0), (-4'h1c), w1, w79, (-31'h14), w97} : {(-6'h10), (-17'h0), (-19'h14), w98, w77, w1, (5'h14), (-32'h1d), w95, (-2'h19), w6, (15'hf), (-22'h4), (-24'h8), w7, (34'hf), (30'h13), (-14'h1d), (-7'h7), (-25'h4), w93, (-26'h1c), (-24'h13)}), (-7'he), (-17'hf), (7'he), $signed(w1)};
assign w66 = (w74 ? w83 : (+(-23'h1b)));
assign w67 = ((w92 || $unsigned(w4)) ? ((~&(w73 ? w92 : w93)) ^ (~&((-23'h3) - {w6, (9'h1c), w5, (16'h6), (14'h12), (22'h15), w3, (20'h19)}))) : (w7 ? w68 : w9));
assign w68 = (20'h17);
assign w69 = (-$unsigned((({w72, (-8'h12), w7, (11'he), w71, (-9'h19), (9'h10), (-7'h0), (7'h19), (27'h12)} ? w1 : $unsigned(w4)) >> (-$signed((22'h5))))));
assign w70 = ($unsigned(w71) <<< ((-21'ha) ? {w77, w80, (14'hd), w86, (24'h7), w2, (10'h13), (24'h12), (-21'h1a), (-9'h14), (25'h5), w96} : ((w99 ? (-5'h5) : (26'h19)) ? w9 : $unsigned((2'h5)))));
assign w71 = (-33'h5);
assign w72 = (w75 <= (-28'h12));
assign w73 = (-4'h12);
assign w74 = ({{w82, w10, (25'ha), (15'h9), (-25'h16), (26'h2), (24'h16), (30'h2), w3, (-28'h1b), (-19'hc), (-27'h2), w77, w8, w82, w8, w6}, (&(25'h16)), {w96, w1, w75, w100, w89, (3'h1d), w3, (16'h15), (29'h11)}, (-5'h5), (-6'h12), $unsigned((-1'hb)), $signed(w90), w75, (w93 & w7), (w81 ? w87 : (-7'h14)), ((12'h18) ? w95 : (27'h19))} >>> w95);
assign w75 = w95;
assign w76 = w97;
assign w77 = (~^$signed(w88));
assign w78 = w5;
assign w79 = w7;
assign w80 = (+($unsigned(((19'h13) === (^~w97))) | (~&$unsigned($signed(w5)))));
assign w81 = (~&(-27'h5));
assign w82 = w95;
assign w83 = (-16'h7);
assign w84 = (w2 ^ ($unsigned(w92) ? (-15'h5) : $unsigned((10'h17))));
assign w85 = $signed({(w10 && (7'h4)), {(-12'h2), w5, (-18'h6), w98, (-28'h1d), (30'hf), (-8'h16), w3, (9'h1c), w92, w5, (25'hb), w86, (-14'h5), w92, (12'hf), (7'h6), (27'hd), (16'h10), w3, (4'h1e)}, (w3 ? (22'h9) : (-20'h6)), (&w92), w6, $unsigned(w6), (w99 ? (8'h19) : (-26'h13))});
assign w86 = (23'h2);
assign w87 = (!((w5 ? w97 : $signed({w99, (27'h8), w100, w8, w96, (29'h1e), w4, (-8'h11), (20'hd), (-30'h8), w94, (-1'h1c), (21'h1e), w97, w3, (20'h6), w6})) <= (+(w10 ? w6 : (|(-11'h1d))))));
assign w88 = {(-9'h1), w95, $unsigned($unsigned((-30'h5))), (+(29'h9)), (w1 ? (w97 || w1) : w96), ((w89 ? w4 : w91) ? (~&(-28'h5)) : (w8 >= w91)), ((~^(19'hf)) ? (+w9) : (-(3'h1e))), (~&{(29'h13), w91, (24'h12), w7, (10'h1c), (-27'he), (6'hc), w4, (-23'ha), (-4'h10), (-8'hb), w92, w3, w97, w96, (19'h16), w93, (-5'he), (15'h2), w92, (-30'h0), (30'h1e), w5}), (-11'h13), ((-21'h18) == ((11'h1b) < (24'h1)))};
assign w89 = (1'h11);
assign w90 = (w2 ? (((11'h15) ? w94 : (w10 - (-9'h13))) ? w10 : ((-24'h18) ? w8 : {(-4'hd), w1, (-6'he), (-21'h0), (-15'h5), (-17'h1e), w1, w5})) : ((-(w4 ? (19'h17) : (12'h3))) !== (-22'he)));
assign w91 = (-22'hb);
assign w92 = {$signed($signed((-16'h18))), ((~&(17'h19)) ~^ ((17'h16) >= w9)), (+(-15'h1d)), ((-2'h9) != $unsigned((11'h6)))};
assign w93 = $unsigned($unsigned((~^$signed({w99, w98, (-12'h0), w1, (8'he), w7}))));
assign w94 = (($signed($signed(w98)) ? ((-11'h17) ? (22'h11) : (w7 ~^ (27'h18))) : ((23'h1e) - ((~^(6'h1)) >>> $unsigned(w98)))) ^ $signed((20'h1c)));
assign w95 = $unsigned(w97);
assign w96 = {(((-6'h19) ? w9 : (-1'h4)) ? w10 : $signed((4'h3))), ((w9 ? w4 : w100) ? ((1'h1d) ? w1 : w98) : {(-25'hb), w97, (4'hf), w8, (-5'h15), w6, (-3'h12), w97, (-16'h1d), w4, (-15'he), w8, (-22'h1c), w3, (4'h1e), w99, (3'h7), (28'h15), w9, (4'hc), w10, (8'h1), (25'h4), (26'hb), (15'h13), w3, (-19'h3), w2, w100, w97}), (+(-18'h2)), (20'h11), (~|w6), {w3, (-18'h7), w10, w100, (1'hb), (6'h15), w6, w2, w3, (5'h16), w6, (15'h13), w100}, (23'hb), (13'ha), $signed((w5 && w98)), (-14'h2), $unsigned(((-5'h7) ? (24'h13) : (12'h7))), w100, $unsigned((~^w7)), w4};
assign w97 = {(~^w8), {(2'h6), (20'hc), (-22'h3), w1, (-26'h1e), w4, w2, (4'h9), (28'ha), (-11'h16), (12'hb), w100, w2}, ((w99 || w5) ? $signed(w4) : ((5'h16) ? (-9'h8) : (30'h1c))), $signed((16'hd)), ((23'h11) - ((-9'h1d) ? w3 : (20'hb))), {(16'h5), w4, (2'hc), w5, (-12'h6), w99, (21'hb), w98, (-10'hf), w8, (15'h15), w3, w8, w8, w10, w10, (11'h2), w9, w10, (-6'h5), (10'h1e), w3, (-25'hb), (-5'h0), w1}, ((w6 * w3) * w7), ((w1 ? w100 : (17'h16)) + (w7 ? (-22'h14) : (-7'h6))), ((~&(21'hb)) > (6'h3)), ($unsigned((-26'h3)) ^~ (24'h3)), w7, {w6, (-26'h12), (20'h1e), (6'hd), w9}, w7, ({(-2'h17), (3'h11), w99} ? {(-22'h12), w6, w10, (-1'he), (21'h5), (-17'h15), (-6'h0), w99, (18'h4), w10, (29'h17), w100, (23'h1b), (16'h1), w3, (2'h17), w5, w8, w7, (-14'h11), w100, (5'h11), (7'h1d), w9, w9, (25'h18), (2'h18)} : (17'h5)), ((5'hd) ? $unsigned(w6) : {w7, (-1'h6), (10'h16), w99, w6, (1'h8), w7, (-5'hf), w3, (-31'hd), (9'h13), (-2'h4), w1, (-24'h3), w2, w99, (-16'h0), w99, (-24'h2), (-13'h4), w3, w4, (-16'h15), w99, (-18'h8), (12'h1c), (8'h3), (-1'hc), (-23'h10)}), (-15'ha), w7, ((-13'hd) ~^ (w6 == (-8'h16))), {w1, (-13'hb), (-18'h17), w2, (29'h1e), w3, w2, w8, w3, w99, (26'hc), w3, (31'h7), (4'h13), (13'h7), w99, (11'h8)}, (w98 ? (~&(-7'h8)) : (-19'hd)), (+(~^w98)), {w100, w98, w3, (7'h12), (-3'h15), w1, w98, w6, w3, w3, w99, w2, (19'h4), (16'h7), (28'he), (11'he), w1, w7, w7, w3, w6, (-16'h1c), (3'h16), (-30'h5), w8, (24'h19), (29'hf), (19'h11), w4}, {w1, w99, w4, w2, w6, w5, (-1'h14), w99, (1'h14), (-14'h1), (3'h9), w99, (-16'h1a), w100, w6, w3, (10'he), w99, (22'hd), w3, (-14'h3), w7, (-4'h1a), (-28'h9), w10, w1}, (|((-9'h1) || w2))};
assign w98 = $unsigned({(5'h4), (w99 * w10), (w4 === w6), (^w5), {(-8'h3), (18'hb), (-15'hd), w6, (-1'h19), (15'h1d), w5, w2, (-7'hf), (29'hd), w5, (29'hf), (-26'h3), (23'he), w8, w8, (16'hc), (-3'h3), (19'h17), w9, (-15'h19), (7'h1e)}, (!w5), ((28'h8) ? (27'h18) : w100), (w1 - (-1'h18)), ((-21'hd) ? (29'h18) : w99), (w4 ^~ w7), (&(-19'h10)), $signed((-24'h19)), (w1 ? (-2'h5) : w10), {w7}, (!(5'he))});
assign w99 = ((-10'h18) ? (|(&((30'h19) ? w8 : (30'h5)))) : (-22'h18));
assign w100 = (-13'h1e);
assign y = {w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100};
endmodule
