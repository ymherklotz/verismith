module test_module(y, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10);
output wire [1505:0] y;
input wire [12:0] w1;
input wire [2:0] w2;
input wire [16:0] w3;
input wire [8:0] w4;
input wire [15:0] w5;
input wire [22:0] w6;
input wire [8:0] w7;
input wire [16:0] w8;
input wire [17:0] w9;
input wire [20:0] w10;
wire [2:0] w11;
wire [15:0] w12;
wire [8:0] w13;
wire [10:0] w14;
wire [28:0] w15;
wire [23:0] w16;
wire w17;
wire [10:0] w18;
wire [8:0] w19;
wire [8:0] w20;
wire [28:0] w21;
wire [10:0] w22;
wire [6:0] w23;
wire [5:0] w24;
wire [22:0] w25;
wire [15:0] w26;
wire [27:0] w27;
wire [18:0] w28;
wire [13:0] w29;
wire [19:0] w30;
wire [1:0] w31;
wire [14:0] w32;
wire [29:0] w33;
wire [25:0] w34;
wire [18:0] w35;
wire [19:0] w36;
wire [17:0] w37;
wire [2:0] w38;
wire [15:0] w39;
wire [21:0] w40;
wire [27:0] w41;
wire [23:0] w42;
wire [14:0] w43;
wire [28:0] w44;
wire [10:0] w45;
wire [15:0] w46;
wire [17:0] w47;
wire [4:0] w48;
wire [26:0] w49;
wire [27:0] w50;
wire [21:0] w51;
wire [23:0] w52;
wire [5:0] w53;
wire [12:0] w54;
wire [15:0] w55;
wire [25:0] w56;
wire [26:0] w57;
wire w58;
wire [14:0] w59;
wire [19:0] w60;
wire [28:0] w61;
wire [10:0] w62;
wire [11:0] w63;
wire [19:0] w64;
wire [17:0] w65;
wire [1:0] w66;
wire [21:0] w67;
wire [14:0] w68;
wire [5:0] w69;
wire [18:0] w70;
wire [26:0] w71;
wire [26:0] w72;
wire [2:0] w73;
wire [2:0] w74;
wire [15:0] w75;
wire [10:0] w76;
wire [19:0] w77;
wire [16:0] w78;
wire [9:0] w79;
wire [8:0] w80;
wire [8:0] w81;
wire [24:0] w82;
wire [28:0] w83;
wire [10:0] w84;
wire [29:0] w85;
wire [18:0] w86;
wire [6:0] w87;
wire [18:0] w88;
wire [27:0] w89;
wire [24:0] w90;
wire [11:0] w91;
wire [13:0] w92;
wire [9:0] w93;
wire [16:0] w94;
wire [25:0] w95;
wire [16:0] w96;
wire [21:0] w97;
wire [18:0] w98;
wire [25:0] w99;
wire [6:0] w100;
assign w11 = (^{(w10 ? w30 : (26'hb)), (w89 ^ w59), (-2'h19), (|(-19'h6)), w93, ((13'hf) ? w20 : (11'h17)), {w15, (1'h3), (-29'h1c), w64}, (w87 && (-6'h13)), (^w85), $unsigned(w21), (~^(17'h1e)), (w3 ^~ (-22'h19)), $unsigned((-29'h15)), (-(-19'h7)), (w40 <= (-22'h17)), ((-29'h6) ? w41 : (-16'h17)), {w78, (-25'he), (30'h1), w1, (-12'h9), w13, w81, (-30'h15), (8'h1c), w73, (17'h1), (-17'h1b), (30'h9), w68, (12'h1d), w12, w42, (-6'h17), w73, (10'h1b), w10, (-8'h12), w28, w74, (24'h10), (30'h17), (2'h1c)}, (w13 ? w81 : w12), {(-7'hd), (2'h5), (-25'h1e), (6'h4), (20'h11), w3, (14'he), (21'h15), (-2'h1d), (14'hc), (-24'h1), w40}, {w49, (-23'h2), (23'h7), w67, w39, (-29'hb), w61, w18, (-24'ha), w93, w37}, w39, ((8'h16) >= (18'h1c)), (!(-3'h16)), (~|(-22'h1a)), {w92, (25'h15)}, {w98, w43, (-26'h1), (-1'h16), (-23'h1d), (-18'h1b), w5, (14'h1), w26}});
assign w12 = ((({(-7'h4), (10'h10), (3'hc), (26'hf), (-18'h1), (-22'h1e), (27'h8), w84, w60, (22'h8), w4, w65, w92, (-30'h17), w10, (16'hc)} ? (6'h17) : (|(w40 ? (23'h19) : w67))) ^ (w90 ? (-18'hd) : ((-12'hb) ? w81 : w54))) >>> w65);
assign w13 = (w64 ? (-15'h14) : (~&(~|{w9, w83, w68, (-11'h12), (-6'hb), w96, (25'hd), (-12'h0), w62, (-5'h18), w44, w41, (8'h1e), (-4'h1), w44, (-30'h1d), (16'h1c), (3'h14)})));
assign w14 = w50;
assign w15 = {(^~$unsigned(w21)), ($unsigned((11'h16)) - (~&w24)), {(31'h4), (-35'hc), (1'h1d)}, ((^(-25'hf)) ? (24'h1e) : (w67 ? w81 : w84)), {(-20'h14), (-25'hf), (-17'h5), w54, (2'h13), (-29'h5), w37, (-10'ha), w70, (-16'ha), (14'h1e), w56, w67, w82, (17'h14), (20'h1)}, $signed((-15'hd)), (~^{w87, w74, w35, w47, (-31'h17), w70, (3'h3), w64, (-5'ha), w44, w41, w76, w47, (-18'h15)}), $unsigned((w70 - w31)), {w34, (-12'h1b), (-5'h1d), w20, w33, w4, (17'h1b), w4, (-13'h17), w48, w25, w48, (-10'h17), w25}, (-11'h8), $signed((w96 ? (-9'h1e) : w38)), $signed((^~(-19'h3))), ((!w30) === (~|w24)), (^~(24'h14)), (+(^w100)), (~&w67), (-19'h0), (-3'h7), (14'h9), ((-(22'ha)) <<< w55), w6, {(-12'hb), w51, (20'h6), (-5'h1b), w4, w25, (-15'h1a), w17, (3'h10), w68, w45, (-4'h1e), (-5'h19), (-13'h12), w75, (9'h1a)}, (-13'h0), ((-8'h8) ? {(23'h18), (-9'h18), w81, w20, w4} : {w51, (-25'h12), w70, (18'ha), w23, w80, w48, w41, (11'h1e), w35, (9'ha), (14'hf), w44, (12'h3), (12'h2), (13'h7), w82, w18, (7'h1b), w62, w58, (7'h2), w2, w31, (-21'hc)}), (w5 ? (w56 ? w56 : w24) : (7'h1a)), (-22'h5), (17'h19), w45, {w53, w98, (12'h14), (25'he), w92, (-9'h1a), w79, w28, (-28'h2), (29'h1b), (-23'h8), (27'hd), w19, (2'h3), w32, w65, (-25'h5), (-23'h16), (-19'hb), (14'h6), w39, (14'h14), (3'h12), (-20'h9), w66, w24}, {(-3'h14), (26'h10), (-10'h16), (-20'h19), (-21'h1c), w83, w23, w40}};
assign w16 = (-15'h15);
assign w17 = ($signed(((!(w89 ? w96 : w46)) ? $unsigned($unsigned(w81)) : {(16'h14), w40, w95, (-9'ha), (4'h1d), w7, (-24'h10), (-6'h15), w36, (-4'h10), (-3'h1c), w73, w83, w34, (-26'hf)})) > ({(6'h7), w33, w83, (1'h1), w47, (-17'hf), w9, w20, (-6'h7), w10, w64, w20, w20, w60, w4, w2} | (-9'hd)));
assign w18 = {(|((-23'h1d) ~^ w23)), {w94, (2'h5), (-14'h18), w96, (-28'h18), (3'h2), w31}, w26, (-(17'he)), (-4'h16), $unsigned((-31'h1b)), w96, (w53 ? $signed(w22) : (20'h1)), $unsigned((15'h1b)), {(-16'ha), (15'he), w79, w9, w91, (22'h18), (-17'h7), (12'he), w53, (-18'hb), w31, (25'h2)}, ($signed((-15'h2)) ? w4 : ((-12'h10) ? (15'h16) : w4)), $signed({w75, (13'h16), w49, w37, (3'h7), w69, w1, w95, (8'h1), (-23'h5), (18'h5), (5'h18), (-20'h3), w72, w63, w74}), $unsigned(((1'h8) != w6)), (((15'h15) ? w76 : (-29'h4)) * (20'h1)), ((w9 ? (-26'h10) : (18'h16)) == (w56 == (16'he)))};
assign w19 = (-{((3'h1b) ~^ w51), (-(11'h7)), $unsigned((-27'h1b)), (w30 ? w48 : w78), $unsigned(w71), {w75, (12'h11), w69, w32, (30'h18)}, (22'h2), w30, $signed(w35), w90, w92, ((-29'h14) ^~ (-26'h1e)), (|w81), w82, (w7 ? w52 : (14'h10))});
assign w20 = {((w97 ? w33 : (2'h2)) ? $unsigned(w26) : ((3'h5) ~^ w57)), (^~(w28 ? (-10'hc) : (26'hf))), ($unsigned((-14'ha)) <<< (~|w39)), (13'h2), (((10'hc) ? (6'h8) : (-1'h1)) < (^(-11'h1b))), (-17'h2), ((w22 <= (23'h16)) ? (w76 ? (11'h16) : (-25'h1d)) : {(12'h4), (25'h15), (-16'h14), w1, (-29'h16), (20'h17), w90, w96, (23'h1d), (3'hd), w94, w67, (-27'h1d), (-21'hc), w57, w73, w71, w10, w96, (23'h6), w85, (32'hd), (-10'h2), (-25'h6), w60, (1'h5)}), {w47, w88, (-5'ha), w99, w100, w81, (-24'h15), w28, (-23'hb), (-17'h6), (-15'h9), (7'ha), w37, w55, (-24'h10)}, ((-22'h13) ^ {(-11'h13), w22, (2'hb), w55, w91, (-27'h6), (-29'hd), w96, (-6'h13), (-27'h16), (22'hb), w33, (-5'hf), w1, (-12'h1a), w83, w35, (-23'h7), w86, (4'h10), w77, w73, w92, w21, w70, w97}), (28'h8), ((w87 | w5) ? w43 : {w99, w36, (-29'h1), w34, w30, (-7'he), (-29'h17), w4, (-5'h13), w62, w6, w28, (-30'h15), (-18'h8), w84, w54, w45, w25, w46, w5, (-10'ha), w29, w40, (15'h1e), (-12'he), (23'hd), w35, w64}), $signed((13'hc))};
assign w21 = ((-7'h12) ? (w71 <<< (&(4'h11))) : (w67 <<< ({w2, w60, w38, (12'h4), (-1'hb), w39, w50, (-1'he), (16'h1a), (-31'h13), w61, (-17'h1b), w34, w29, w22, w68, (8'h3), (1'h1c), (12'h5)} ~^ ((|w38) & ((-2'h12) ? (-18'h8) : w84)))));
assign w22 = ((w61 && ((w44 ? (-11'h19) : (-19'h6)) ? (^(!(-1'h8))) : ((-24'h12) ? (27'h6) : w70))) <<< w84);
assign w23 = w68;
assign w24 = (-8'h3);
assign w25 = (24'ha);
assign w26 = (&{(-14'h3), (12'h8), (10'h19), (25'h17), (w96 - (27'h4)), {(-5'h16), (-26'h6), (-24'h4), (21'h13), w64, w81, w6, w81, (5'h7), (3'h2), (19'h16), (-29'h1c), w2, (29'h3), (-4'h14), w99, (-9'h9), (-12'h15), w53, (14'h1c), w42}, w65, (2'hf), (w5 !== w30), ((-6'h19) ? w95 : (-23'h1a)), $unsigned(w53), (^(22'h9)), (w96 ? w82 : (13'hb)), w35, w9, $signed(w72), (+(10'h1b)), {(-16'h17), w40, w56, (16'hb), w64, (-11'h15), w68, (32'h18), (-14'h13), (6'h4), w82, (-26'h16)}});
assign w27 = (($signed((-17'h2)) & ({w42, (12'h18), (-28'h1c), w7, w92, w8, (10'h2), w97, w2, w57, w97, w71, (1'h4), (16'h13), w47, w89, (4'hf), w72, w32, (-22'h6), w66, w68, (-30'h0), w48, w70, w44, (-3'h15), w63, w76, (26'h5)} ? ((~^(32'hd)) >= {w89, (18'h1d), (5'hb), w57, (-30'h2), w94, (15'h16), w38, w70, (-5'ha), (17'h9), w39, w45, w72, w79, w39, (25'h7), (-8'h13), w30, w29, w51, w59, w7, w82, w92, (3'hf), (-20'h1a), (17'hc), (28'ha), (11'h9)}) : ((-16'h12) ? (23'h16) : (30'h3)))) || (-30'h1));
assign w28 = ((($signed((14'h19)) << (&w30)) ? $signed((!(21'hc))) : (-14'h1e)) ? w80 : {((24'h3) ? (19'h12) : (-7'hf)), (&(9'h13)), ((-3'h16) - (-35'h12)), (w45 ? w94 : (29'h17)), (w45 ? (24'hd) : (28'h17)), (w73 ? (17'hf) : (-29'h13)), $unsigned((-36'h8)), $unsigned(w99), (w91 | (29'h4)), {w73, (17'h2), (-26'h1b), w67, w86, (2'h8), w79, w44, w78, (-9'he), w43, (30'hb), w33, (-8'h19), (-17'h1), (-23'h6), w86, (-8'h19), (12'h16), (9'hd), (10'h15), w49, w35, (-1'h10), (20'h11)}});
assign w29 = (-27'h4);
assign w30 = w60;
assign w31 = (6'ha);
assign w32 = w43;
assign w33 = $signed($signed((-6'hf)));
assign w34 = w78;
assign w35 = $signed({w61, ((-13'h16) ? (-15'ha) : (33'h18)), ((20'h13) ? w75 : w40), w39, ((19'h1c) ^~ (7'ha)), ((16'h17) - (-20'h5)), w36, (~&(17'h17)), w67, (^(10'h11)), ((9'h13) ? w84 : (-25'h16)), (w49 ? (-15'hd) : w79), {(19'hc), w49, (-26'hb), (30'h1c), w92, w68, w72, (17'h3), (5'h14), w99}, ((19'ha) && w63), (&w43), {(11'h10), (-4'h10), (-30'h0), (-28'h15), w38, (3'h2), w99, w39, w85, w63, w79, (22'hc), w48, w99, (14'h16), w56, w40, (27'h1c), (16'hc)}, {w63, (-15'h1a), (-1'h2), (-22'hc), (1'h13), (16'h3), (-18'h1d), w66, w92, w41, w95, w51, w3, w43, (-7'h1e), (6'h1e), (-29'h18), w47, (29'h13), w70, w78, w50, w66, w45, (-26'h2), w53, w92, (22'h5), (-14'hc), w10}, ((3'h4) || (20'h6)), {(7'h18), w86, w84, (-21'h18), (6'h1b), w61, w9, (-7'hf), w73, (17'h1), w96, (-8'h16), w84, w40, w73, w48, w9, w57, w80, w87, w95, (22'h18), (17'h17), w66, w43}});
assign w36 = $signed($signed(w5));
assign w37 = ({(w86 ? w51 : (11'h14)), (^~w87), {(9'h6), (22'h1b), w10, w57, w56, (3'hd)}, w49, ((-34'hd) ? w88 : w3), (-15'h18), (+(-11'h8)), w59, (-5'h7), $signed((-19'h1a)), (w44 * w50), (~&(-28'h1e)), (w43 * w97), ((-8'h1d) ? w89 : (-18'h1b)), $signed(w49)} | {(^~(13'h14)), w74});
assign w38 = (~&(28'hb));
assign w39 = {(11'h16), ((-36'ha) ? (~^(-32'h16)) : ((-13'ha) + (21'h14))), ((w1 && w57) - {(3'h19), (-20'h1a), w85, (-23'h18), w85, w88, w68, w56, w54}), (-{(28'h8), (15'h1a), (10'hd), (-17'h11), w56, w55, (-27'h14), (-7'h12), (-10'h12), (-34'hd), (22'h17), w79, w88, w46, (7'hb), w59, (-26'h12), w6, (26'ha), w88, (27'h1c), (-9'h14), (-15'h11), w70, w87, w3}), {(-32'h1b), (-16'hc), (29'ha), (-24'h5), (-28'h8), (8'h1b), w76, w41, w75, w94, (23'h3), w45, (21'h6), (-26'h1c), w82, w57, (-7'h2), w43, w98, (-18'h18), w56, (-8'h1a), w95, w97, w62, (-8'h8), (24'h3)}, (w82 >> $signed(w88)), {(16'hb), (22'h1e), (5'h7), (-7'h17), w70, w63, (2'ha), (16'h15), w49, (-16'hf), (-9'h1d), w53, (19'hb), (-22'h14), (-13'h18), w66, (-28'h14), (24'h1d), (-28'h1), (-2'he), (11'h1e), (-12'h17), w56, (1'h17), w95, w42, (1'h5), (-19'h0)}, $unsigned(w55), ((&w8) ? w60 : $unsigned(w59)), {w72, (-15'h11), w2, w63, w59, (10'h1a), w48, w71, (-27'hf), (-29'h17), w91, (-8'h1a), (-11'h4), (7'h15), (-26'h15), (10'h16), w7, (-29'h11), w81, (12'h4), (23'h8)}, w56, $unsigned(((1'h2) ? (4'h6) : w98))};
assign w40 = $unsigned({((27'h1a) ? (31'h17) : w92), {(-31'h1), (-10'h7), w9, w83, w2}, (w78 ? (-7'h2) : (-2'h1b)), (28'h13), (23'h3), (-16'hc), (|w46), $unsigned((-23'h1c)), (w50 ? w72 : w100), (6'hc), (w87 ~^ (-26'h1a)), (w89 >= w88), (30'h8), w87, $unsigned((21'h8)), (^(12'h1c)), $unsigned(w96), (-15'hb)});
assign w41 = (20'h19);
assign w42 = ($unsigned(w97) ~^ $unsigned((19'h1c)));
assign w43 = (-27'h10);
assign w44 = (-29'h19);
assign w45 = {($signed(w46) ? ((24'h10) << w93) : $signed(w78)), ($unsigned(w93) >> (~&w84)), (^((-21'h16) >= (29'h11)))};
assign w46 = {$unsigned(w68), (&(20'h18)), w98, (-9'h1c), {w72, w47, w74, w88, (-25'h3), w62, (12'h15), (29'h9), w80, w66, w63, w70, w67, (16'h4), w70, w1, (-6'hb), w56, (-26'hb), (25'h1b), (24'hb), (-20'h11), (13'h5), (-5'h7), (-6'hf), (-21'h1d), (-7'hb), (-28'hb)}, ({(-17'h1e), (-12'h1d), w5, w92, (22'h1a), (6'h15), (18'h12), w77, w97, w58, w64, (6'h2), (-27'h2), w47, w9, w81, (18'hd), (9'hc), w97, w57, w96} >>> w76), $signed({(11'h5), w53, (8'h1e), w99, w100, w83, w62, w68, w79, w83, w62, (31'h1c), (15'h3), w77, (1'h11), (6'h19), w8, w63, (-23'h9), (10'h15), (-26'h18), (-25'h1d), w59, w99, w89, w64, (13'h1b), w50, w98, w76}), $unsigned($signed(w74)), $signed((-31'h19)), ({w97, (26'h1), (20'h15), w50} ? ((-21'hf) ? w63 : w83) : (16'h10)), {(25'hd), w94, (22'hb), w78, (1'h12), (12'h1b), w91, w5, (-8'ha), w47, (9'h1e), w49, (-32'hf), (-11'h7), w76, (6'hb), (2'h1a), w68, (-20'h6), w58, (-16'h1b), w79, w1, w81, w62, w75, w85}};
assign w47 = ((5'h10) ? ($signed((&(-16'hd))) ? (27'h19) : w78) : {(-5'h15), (w88 ? (-19'hb) : (-19'h0)), $unsigned((14'h3)), $unsigned((-23'h10)), $unsigned((-25'h7)), w54, (-(11'h11)), ((1'h9) && w96), (-10'h5), $unsigned(w95), {(30'h16), (-19'h10), (-27'hd), (17'h1e), w69, (-5'h7), (-29'h13), w66, (-8'h9), (-9'h15), w94, w76, (-20'h16), (4'h2)}, ((-17'h16) <= w75), w53, $unsigned(w58), {w89, w68, w88, (-28'h17), w53, (20'h3), (7'h4), w76, (8'h17), w55, w1, w67, (18'h1b), w82, w10, w98, w70, (-23'h15), (12'h1e), w64, (20'h10), w63, w5, w60, w81, (11'h13), w76, (8'h17), (-1'h14), w68}, w94, w93, (+(19'h13)), $signed((6'h2)), {w78, w61, w65, (-28'h17), w54, (27'h8), (-21'h4), w72, w1, w83, w66, (-7'he), w93, (-13'h3), (4'hf), (-12'ha), w55, (-22'h3), w54, (-10'hc), w55, (11'h1e)}});
assign w48 = {(-(11'h9)), {(-29'h4), (23'h17)}, ((^(17'h8)) ? (|w57) : {w10, (-32'h14), w64, (-20'h19), (5'h1b), w7, (17'h17), (12'h10), w65, (16'h13), w51, (-5'ha), (-14'hd), w10, w53, (30'he), (27'h19), w53, w71, w90, (19'h9), w86, w8, w72, (-9'h12), w71, w73, (16'he), (-29'he)}), {(10'ha), (-18'h4), (-22'h14), (20'ha), w61, w68, (19'h16), w4}, (~|$signed((11'h12))), (((19'hd) ^~ (-19'h0)) ? (+w66) : w99), {(-21'h1c), w65, (-15'h16), (-32'h5), (29'h16), (-8'h14), (8'ha), (19'h3), w6, (25'h17), w72, w70, w4, w72, w60, w88, w77, (13'h18), w3, w63, w98, w96}, w86};
assign w49 = (-10'h1b);
assign w50 = $signed(({w89, w86, (22'h8), w81, (25'h3), w59, w78, (-15'h14)} >> $unsigned($unsigned((~&w78)))));
assign w51 = $unsigned({(24'hf), (!(13'h16))});
assign w52 = (-7'h15);
assign w53 = (({w8, (-11'h1), (-28'h1a), w64, (1'h1a), (8'h12), (21'h17), w98, (-21'h17), w78, (3'h1d), (24'h18), (-1'ha), (13'h1), (28'h18), (18'h4), (-11'h18), (-9'h8), (-10'h16), (-14'h5), w74, w92, w81, w59} ^ (~&(-7'h1))) < $signed((-7'h1a)));
assign w54 = (^((((w73 <= (11'h7)) > (^~w9)) ? ((18'hb) ? (-14'ha) : (-15'h9)) : $signed({(17'h1b), (16'ha), w84, w82})) <= w79));
assign w55 = ((-28'hc) ? w62 : ((|(~&w67)) ? (-((8'ha) ? (-32'h3) : (-17'h19))) : $signed(((-7'h7) ? (23'h8) : w59))));
assign w56 = (~&w68);
assign w57 = ({(25'h5), w79} + (w87 ? w76 : (-8'h10)));
assign w58 = ({w74, (w92 ? w6 : (-27'hf)), ((5'h1b) ? (18'h1d) : (-9'h1c)), (~&w59), (w82 ? (30'h4) : (6'h16)), (~&(30'hf)), (w77 ~^ (20'hf)), (!w92), (19'h3), {(-8'h1e), (25'h17), (19'h4), (-16'h9), (-16'h1a), w86, w9, w63, (-19'h6), w80, (-5'hb), (-29'h11), w80, (-5'h17), w98, w84, (17'h9)}, (w96 ^~ (2'he)), (-1'h18), (30'h12), (-13'h1a), w5, {w79, w59, w6, (3'h10), (-15'h16), (-23'h5), (17'h1e), (25'h12), w86, w92, w85, w72, (-20'h0), (-24'h3), w94, w65, w88, (-12'h2), (-14'ha), (30'h1a), w68, (7'h1a), (-2'h19)}, w78, ((18'hf) ^~ w67), (~|(26'h1a)), (-14'hd), $unsigned((-6'h1c)), {w65, (29'h19), (18'hf), (-26'hf), w97, (-19'hf), (26'h1), (28'h10), w72, w81, (19'h19), w60, w87, (-26'h16), (-7'h9), w73, (-31'h19)}} > (|(((15'h3) ? (2'h19) : (16'h19)) ? w10 : (&{(6'ha), w62, w73, w83, (-9'h2), (-17'h1c), (11'hf), (-28'h12), (-27'h8)}))));
assign w59 = {{(-33'h1c), w68, (5'h1d), (-10'h4), (-13'h1b), w5, w75}, w97, (^(15'hc)), ({(-20'h13), (16'h4), (21'h1c), w8, w82, w62, (-11'h1), w95, (-26'h3), w6, (-5'h1c), (-20'h10), (7'h1d), w6, (-9'hf), (26'hc), (13'h3), (24'h10), (3'h5), (10'hd), (-8'h1b), (-5'h4), w2} ? w98 : (w90 | (-4'h16))), w5, (3'h1), w85, (~&w67), w76, ($signed(w68) || (w95 ? (-12'hf) : w84)), {w3, (23'h1c), w86, (-21'h18), w97, w10, (-15'h4), w4, (30'hc), w65, (-10'ha), w63, (19'hb), (31'h8), w61, (6'h19), (10'hc), w8, w90}, (&((9'h1a) >= (27'h6))), ((~&w87) != ((11'h4) ~^ (13'h16))), w1, (w3 < ((16'h13) !== w66)), (-{(4'h1c), (-14'h2), w6, (12'h1e), (-21'h3), w68, w71, w88, (-2'h8), w4, w96, (28'h12), w63, w8, w72, (1'hb), w2, w98, (14'h8), w83, (-1'h1d), w75, w71, (-1'h5), (-28'hd), w89, w88, w65, w100}), (((-29'ha) ? w73 : w69) ? $unsigned((-11'h12)) : $signed((21'h16))), ({w91, w8, w96, (14'h4), (6'h3)} == {(29'h13), (8'h14), w5, (23'h12), w61, (11'h14), w64, w80, (-25'h12), (-2'h13), w7, (-17'h18), w85, (23'h5), (20'h6), w86, (24'h5), w74, (-15'h19), w65, w99, (2'hb), (-9'hb), w88, (-11'hb)}), (^(w7 >= w70)), ($signed((-20'h4)) ? w76 : (w6 ? w2 : (-24'h2))), (w78 ? ((24'h4) ~^ (-25'h1c)) : $unsigned((22'h6))), {(-26'h5), w71, (4'h7), (2'h12), w89, w67, w97, w71, (24'h19), (-12'h1d), w99, (-27'h18), (-10'h14), w75, (23'h1a), w96, w67}, ((-16'h2) ? (w9 ? (-24'h8) : w63) : {w91, w96, (9'hd), w92, (-11'h8), w100, (15'h18), w89, (9'h10), (-32'h17), w9, w61, w62, (16'h4), w100, w95}), ({(16'h10), (-20'h19), w82, (2'h9), w88, (-9'h17), (-6'h16), (-2'h1d), w92, (12'ha), (24'h9), (-16'h5), w9, (18'h9), w72, (-6'h1d), w10} <<< (w7 ? w1 : w80)), (w62 ? (!(-30'hd)) : (w99 <= (30'h1b))), (|(|(-25'h1d))), ((-5'h10) != ((-20'h14) === w75)), {w9, w98, (33'h6), w62, w8, w79, (19'h1), w6, (6'he), (-1'h2), w95, (4'h15), (26'h1), (2'h2), w63}};
assign w60 = {w78, w79, ((w90 ? (-7'h1) : (20'ha)) || (-23'h10)), (^~(-11'h1e)), ({w82, (-1'h17), w91, w3, (2'h1a), (21'h19), (14'h12), (31'h14), (-10'h0), w2, (-33'h11), w7} && w81), (w96 <= {w88, (14'hc)}), w81, (-7'h1c), ($signed((-15'h16)) + (~^(-9'h1c)))};
assign w61 = $unsigned(({w100, w64, (-12'h1), w96, (-13'h15), (22'ha), (-29'h9), w2, w9, w2, (8'h16), (26'h19), w93, w7, w88, w69, w67, w95, (-29'h15), w5} ? w65 : ((w74 !== (16'h1)) ? ((-27'h16) >= w85) : (18'hc))));
assign w62 = ((&(4'h11)) + $signed((w84 ? (10'hc) : ($signed((-20'ha)) <= (w8 ^~ w86)))));
assign w63 = w67;
assign w64 = ({(15'hf), (-10'hc), ((18'he) !== w84), ((6'h15) ? (-3'h0) : (9'h1d)), (w10 ? w84 : w93), {w93, w66, (2'h16), (2'hb), w98, w2, w9, (-19'h13), w2, w2, (-22'h13), w80, (-14'h4), w2, (16'h12), (11'he), w84, (-8'h3), (6'h9), w71, w91, w65, (-23'h16), w1, (-2'h17), (-30'ha), (-30'h17)}, (w87 ? w78 : (-2'h11)), (!w94), {(9'h1d), w2, (12'h17), (24'h8), (21'h14), (21'ha), (9'h2), (8'h13), w85, w87, w65, (23'h2), (17'hf), (8'h3), (11'h14), w82, (-28'h1), w1, (-29'h7), w9, w9, (5'h17), w98, (29'h1b), (6'h19), (27'h5), (16'h13), (-29'ha), (-20'h1e), w94}, (~&w100), w91, (^w73), (w78 ^~ w69), (26'h1b), $unsigned(w5), (w74 ? (-20'h18) : (-2'hf)), (23'hb), (-26'h1b), ((-3'h14) - (26'h10))} >= ((~&w94) ~^ $signed(((-31'h2) == w90))));
assign w65 = $signed(((24'h1) ? w67 : {(-4'hb), w9, w82, (9'h1), (-18'h13), w81, (-21'h17), (2'hb), (-10'h1c), (-13'h4), (-21'h1d), (-11'h15), w8, w72, (-23'h13), w10, w67, w97, (3'h10), (-9'h7), (-19'h13), (35'h1b), (19'h5), w6, w3, w67, (28'h1e), w86}));
assign w66 = {(^((18'ha) <<< w68)), $unsigned({w86, (-4'h15), (14'h13), (-6'h1c), (5'h1e), (31'h15), (-15'h1d), w80, w9, w8, w93, (-30'hc), w76, w89, w97, w88, w5, (33'h1d), w87, w84}), (^~(-2'h18)), (~|{w71, w93, w90, w7, (7'h15), (-23'h8), (-27'h2), (26'h6)}), (29'h1a), w89, (4'h1b)};
assign w67 = (-14'h2);
assign w68 = w82;
assign w69 = (w5 ^~ {((12'h1d) ? w96 : w3), {(26'hd), w3, w71, w70, (17'h1c), (18'h15), (-27'hf), (16'h10), (-25'hb), (-25'h11), (-27'h0), w99, (-9'h17), w89, w88, (-13'h1d), (-6'h1a), w79, (6'hf), (3'h19), (-23'h5), (25'h1a), w90, w2, w3, (26'he), w89}, (^~w1), (w79 ? (25'h3) : w4), $unsigned((-6'h16)), ((10'h19) === w78), (~^(2'h16)), ((-25'ha) ? (25'h12) : (-29'h7)), (w99 ~^ w72), (w71 ? w76 : w81), (w83 ? w84 : w2), w86, (20'h19), (-11'hf), (-22'hf), (w72 ? w100 : (-12'h1b)), {(13'h13), (-25'h1e), w86, w75, (-9'h16), w77, (-5'hf), (-17'h2), w2, w89, w98, (20'h19), w79, (-15'h2), (22'h1e), w82, w81, (-16'h1e), w87, (-18'h0), w2, (14'h1e)}, w77, ((-13'h10) ? w2 : (8'h18)), (-4'h7), w98, (~|w86), $signed(w100), {(24'hc), (-31'he), (12'h16), w10, w86, (-17'h18), w89, w3, w75, (-26'h8), (-21'hb), (-31'h11), (-9'h1a), (29'h13), (30'h14), w100}});
assign w70 = w81;
assign w71 = $unsigned((-17'h11));
assign w72 = ((-3'h13) ? ((-21'h1c) ^ $unsigned((-{(-20'h1b), (20'h13), (4'hc), (-12'h11), w10, (23'h7), w77, (-30'h7), (-2'h4), (-15'h1b), w1, (-7'h5), w81, w89, w81, w97, w94, (14'h2), (-7'h5), w4, (30'h16), (-15'h7), (-17'h8), w4, w97, (32'h1a), (24'h1), w80}))) : (^~$signed((((2'hc) ? w78 : w91) ~^ w7))));
assign w73 = ({{(30'h17), (-27'hb), w97}, (w4 !== (33'h16)), ((-26'hd) ? w92 : (26'h10)), (21'h1), ((-11'h16) ? w100 : w82), (w95 ? w10 : w81), (21'h1b), w89, {(-18'h10), (-18'h1a), (-7'h16), w77, (22'h7), w83, w2, w90, w97, (-19'h0), (-1'h6), w90, w75, (19'h1c), (-22'h1e), w6, w93, w93}, {(26'h16), (-16'ha), (-16'h12), w3, w1, w99, w96, (-16'h10), w95, w5, (27'hb), (13'h2), (17'h7), w84, (9'h12), (-19'h14), (17'h7), w78, (-26'he), w8, w83, w7, w90, (20'h11), w91, w76}, (^~(4'hf))} ? (-3'ha) : {{(-9'h15), w80, (16'h1a), w87, w90, (5'h2), (-12'h14), w78, (2'h12), w78, (-24'h8), w87, w89, w90, w76}, (-14'hc), w86, (~|(-3'he)), w86, ((-2'h16) == w4), (~&w89), (^w78), $signed(w93), ((-10'h17) != w76), (-9'h8), (-(28'he))});
assign w74 = {w80, (6'h4), {(20'ha), (-27'hb), (5'h14), w76, w9, w100, (23'h9), w10, w82, w4, w85, w86, (28'ha), w87, w82, w3, w78, w99, w84, w100, w99, w90, (-27'h10), w1, w93}, (-20'h16), w94, ({w87, (-24'h3), w100, (26'h13), (29'h8), (11'hf), (-5'h1b), w98, w93, (-9'h6), w93, w4, w90, (-22'he), (26'h1a), w91, w2, (24'h17), w95, w85, w77, (5'h1d), (16'ha), (26'h9), (19'h10), w94, w4} ? (!w75) : $unsigned(w87)), w6, $unsigned((6'h10)), $signed({(4'h4), (-22'h2), (27'h16), w10, w2, w98, w1, (-32'h14), (28'hf), (22'h15), w9, w84, (-1'h19), w98, (14'hf), (-28'h4), w94, (31'h3), (-28'h1d), w95, (18'h2), w1, (6'h17)}), w98, w95, (^((5'h16) + w89)), (10'h1e), ((w4 <= w87) ? (!w82) : ((6'h8) >= (-20'hf))), (&w1), {(24'h16), (30'h7), (9'hb), (-15'he)}};
assign w75 = ($unsigned(($unsigned(w3) ? (w76 <= w89) : {w77, (-7'h18), (-14'hc), w86, w79, (26'h1e), w5, (-22'h9), (-25'h1b), (-6'h13), w87, w92, w8, w85, (-3'hb), w78, (-15'he), (31'h15), w8, (11'h3), (4'h19)})) ? $signed(((10'h17) <= ((w93 ? w1 : w7) <<< (-27'hc)))) : {$unsigned((10'h12)), (-(23'h11)), ((-16'h17) ? (5'h9) : (-12'h4)), $unsigned((21'h15)), (w86 << (-13'h13)), (w93 ? w2 : (-28'h16)), (w97 & w92), (~&(9'h1c)), ((26'h1) ? (-25'h7) : (-25'hd)), {w84, w94, (28'h3), w96, (10'h19), w93, (-28'h12), (23'h8), (-9'h0), w76, (-32'h1e), w94, (-6'h14), (-9'h12), w97, w98, w7, w91, w92}, $unsigned(w6), {w76}, (-6'ha), w99, (&w4), {(-30'h1c), (-28'hd), (-27'h15), (-8'h0), w87, (30'ha), w79, w92}, w89, ((30'h5) ? (1'he) : (18'h6)), $unsigned((9'h8)), {w84}, (~|(-25'h0))});
assign w76 = {(13'h15), {w100, (8'h1), (16'h13), (-20'h12), (-2'h8), (24'hc), w85, w1, w6, w81, w99, (31'h7), (4'h6), (-4'h2), w5}, (&(^(-7'h9))), (~&{w94, (15'h17), w9, w93, w3, (2'h1e)}), w91, $signed((w87 ? w9 : w9)), w97, $signed((-21'hb)), (^~(-21'h12)), (^(-24'h8)), {(-30'h13), (-17'ha), (-31'hf), w85, w2, w99, w96, w99}, (w94 !== $unsigned(w6)), (5'h2), ((5'h2) ? ((-5'hd) ? (-14'hb) : w81) : (23'hb)), ((w81 ? (-18'h2) : w91) || (w95 | (-1'h16))), ({w3, w8, (-11'h6), w3, (15'h5), (24'h10), (-9'h18), w83, (8'h3), w82, w81, w78, w83, (-8'h7), w4, (-23'h2), w82, (-17'h11), (-14'h16), (28'h1d), w85, (5'h10), (-7'he), (14'h1e)} || {w99, (-14'h8), w78, w90, w88, (24'h1a), (29'he), (5'hd), (18'h1d), w96, w90, w1, w91, (22'he), (-27'hd), w87, w91, w78, (-10'hf), (-1'h1), w10, (26'h6)}), (((-15'h18) ? (21'h11) : w8) <= (w83 ^~ (-26'h9))), $unsigned({(-13'h5), (-7'h1a), w4, w96, w90, w2, (28'hd), w4, w87, w2, w2, (26'h14), w80, w96, w95, (5'hf), w99, (-25'hd)}), (-21'h6), (w96 ^ (-w9)), w94};
assign w77 = (-7'h3);
assign w78 = w84;
assign w79 = (32'h13);
assign w80 = (-10'h2);
assign w81 = (((29'h1d) !== {w91, (-23'hc), w88, (-3'h11), (-28'he), (3'hf), w85, w2, (26'h8), (-25'h15), w10, w96, (-3'h17), w99, w84, w91, w8, w1, w97, w86, (31'h1a)}) ? (|$signed((14'h12))) : ({(1'he), w3, (11'h19), w88, w9, w2, (27'hf)} ? ((-7'h18) || (27'h9)) : ((-19'h9) - (-25'h1b))));
assign w82 = {{w91, w7, w7, w97, (15'h19), w87, w4, w97, (-25'h0), w8, (3'h4), (-19'he), (33'he), (26'h12), (-20'h1b), (17'h1e), (-10'h1a), w91, w92, (21'h1), (-27'h1d), (-23'h7), w7, w88, w96, (8'h3)}, ((~|(-2'h6)) ? ((19'he) ? (19'h7) : (2'h11)) : {(18'h17), (5'h4), (-21'ha), w1, w7, (13'hc), (13'h1c), (22'h1), (-21'h17), (-31'h3), (25'h6), (-24'h1b), (17'h12), (29'ha), w84, w91, (-16'h4)}), $signed((14'h19)), {w86, w89, (22'h14), w85, w98, w8, w1, w88, w90, (-7'h10), w93, (24'h9), (-21'h1b), w92, (18'hc), (-29'h9), w96, w95, (-14'h6), (27'h3), (-30'h1a), w97, (15'h7), w96, w98, w89, w85, w85, (29'hb)}, {(-9'h19), (9'h9), w88, (-14'h1c), (-9'h1b), (-12'hf), w2, (-14'h3), (6'hc)}, ((5'h1d) ? ((15'he) < w6) : (w6 ~^ w9)), ($signed((9'h6)) == w3), ({w93, (3'h6), w89, (20'h18), w6, w3, w9, w88, (1'h19), (-7'h2), w84, (-4'h5), (-28'h2), w99, w97} > ((6'h10) - w9)), ($unsigned((29'ha)) ? $signed(w9) : {(2'h5), w93, w2, w86, w94}), w1, (11'h10), (!(^~(-17'h6))), {(-14'h1), w89, (27'h15), w4, (-12'h13), w2, (24'h19), (-18'h7), w91, w2, (-19'h1a), (-31'h1c), w86, w1, w96, w9, (16'h3), w86, (11'hc), w83, (-19'h17), w97, w3, w2, (22'hc), (-7'he), (27'h1b)}, (-22'h5), (-10'h3), w8, $signed(w88), ({(-20'hf), (34'hf), (28'h1c), w10, w93, w97, w87, w87, (-12'h4), (-14'h17), (-3'h8), w2, w98} == (w96 ? (16'h2) : (-12'h1d))), (((26'h14) !== w97) << ((26'h1d) ? w95 : w10)), $unsigned((-27'h16)), (!(10'h6)), (+w7), ((5'h17) ^~ w88)};
assign w83 = (-22'h1b);
assign w84 = {{w2, w9, w85, w93, w92, w3, w2, (2'hf), (-8'h8), w94, (-10'h4), (-29'h11), (4'h13), w91, (28'hc), w93, w94, (-12'h1e)}, ((&(-3'h14)) ? (-9'h1) : (!(-6'h1c))), w8, $unsigned((9'h6)), {w87, (16'h5), (-30'h18), w10, (-25'he), w9, (-15'h15), w9, w1, (-11'h19), (-21'h1c), w7, (-13'hc), (2'h12), (14'hc), w90, w85, w96, w2}, $unsigned((~|(-27'h12))), (-29'h13), w96, {(-25'h9), w96, (-27'he), (-19'h5), (-12'h2), (-5'h19), w99, w6, w3, (12'h18), (6'h17), (-17'hb), w89, (1'h2), (-21'h4), (-30'h1e), (-13'he), (29'hf), (5'h13), w7, (-7'h1b), w89, w98, w7, w6, w100}, w95, (-8'hb), (20'h2), $unsigned(((-3'hb) ? (2'hc) : w88)), ((|w86) ? (-(25'hc)) : $signed(w95)), ({(20'h8), w6, w8, w1, w4, (-9'h1c), w94, (21'h11), (-30'h17), (-2'h1d), (27'h6), (-5'h13), (-17'h18), w87, w88, (-29'h1e), (-34'h17), (-4'h6), (21'h1c)} ^ (w96 ? w100 : w90)), {w88, (-14'hd), w88, (10'h9), (-29'h1a), (-15'h9), (10'h13), (5'h2), (28'ha), (15'hf), w97, w91, (-3'hd), (24'hf), (1'h4), w4, w99, (-28'ha), (26'h7)}, w10, ((w4 ? w4 : (-21'hb)) ? (-(-16'h17)) : {w97, (7'hf), (26'hd)}), (^~{w90, w6, (-26'h5), (28'h11), w4, w1, w88, w10, (4'h1c)}), (-w9), (-18'h13), $signed((|w9)), (((7'h1e) == w88) ? $unsigned((19'h11)) : $unsigned((28'h1))), ($unsigned(w93) | {(-26'h1), w3, (5'h15), w92, (25'h3), (-17'h3), (-26'h4), w95, (3'h3)}), (!{(-9'h9), (28'h7), w94, w89, (22'h17), (-26'h18), w86, w89, w4, w9, (17'h6), (-21'h19), (-9'h17), w9, (-4'h1a), w2}), (-31'h1c), ((w2 ? (29'h16) : w98) ? w95 : $signed((12'h17))), ((w97 ? (-3'h3) : w7) - ((19'h1) == w93)), {w86, (-22'h10), w86, w88, (-19'h2), (22'h15), (18'h14), w9, w88, (-2'h6), (-10'h18), w10, (30'h4)}, w100};
assign w85 = {(!w89), ((w99 ? (-12'h1b) : w93) ? $unsigned((8'h5)) : w88), $signed({w87, w98, w97, (-29'h9), (-10'hd), (-9'h10), (-18'h4), (7'hc), (10'h6), (13'h7), (12'h8), w97, (-1'h18), w95, w96, w88, (7'h1b), (-4'h18), w86, w92, (3'h1), w90, w93, (9'h1d), (23'h17), (-9'h17), w91, (3'h8)}), (25'h1c), (~|$signed(w89)), $unsigned((-23'h1c)), ((w5 ? w88 : (14'h12)) ? (w90 < (-30'h0)) : {w89, w89, (2'hb), w1, (1'h1), (16'h1c), w10, w2, (2'h1a), w91, w10, (23'h1d), (18'h16), (-5'h12), w91, w89, (1'h6), (-23'h16), w1, w95, w91, (-8'h0), w9}), $signed((~|w92))};
assign w86 = (15'h14);
assign w87 = ({$signed((-30'h5)), {(-1'h16), w8, w88, w1, w98, w99, (24'h4), (-17'h1e), (-20'h10), (-11'h16), (31'h1b), (-20'he), (3'hc)}, (w94 ? (-4'h1c) : (1'h14)), (^w95), $unsigned((-24'h1d)), w98, (w1 ? (23'hf) : (26'h3)), ((-21'h13) ? w93 : w9), $signed((21'he)), {w98, w4, w98}, (10'h9), (w10 ? (10'he) : w88), {(23'h10), (-29'h17), (15'h12), (21'h1), w93, (15'h1a), (20'h4), (-21'hc), w91, w96, (30'ha)}, (-23'h1c)} + $signed((&(!((-10'h18) * (-13'h1))))));
assign w88 = (($unsigned((-27'h14)) >>> $signed((-$signed(w94)))) - $signed(w6));
assign w89 = $unsigned((11'h13));
assign w90 = $unsigned((~|(&(-26'he))));
assign w91 = $signed(($unsigned((^~(-13'h13))) ? ((w94 ? (-27'h5) : w10) != {(-5'hc), w94, (21'he), w95, (-4'ha), (3'h8), (-30'h1), w1, (-15'h1b), (22'h5), w8, w2, w100, w97, (17'hc), (18'he), (27'h1b), (-17'h1d), w2, (-24'h1d), (22'h13), (23'h14), (15'h19), w1, (13'h15), (10'h3)}) : (19'h4)));
assign w92 = ($unsigned((+$unsigned((w3 & w99)))) ? {(-12'h14), (^w5), ((-8'h8) ? (1'h8) : (11'h7)), (w1 ? (-17'h18) : (-31'h5)), ((-9'h12) ? w7 : w8)} : {(~&w6), (w8 === (-27'h2)), {w2, (25'h15), (6'h1e), (-8'h3), (-6'h17), (-1'h5), (-30'hf), w98, w1, w4, w100, (6'h12), (22'h12), (-26'h11), (-7'h7), w94, (4'h1d), (23'hb)}, (-w10), $signed((14'h1)), w99});
assign w93 = (-24'ha);
assign w94 = {w4, (((26'h9) ? (2'h1a) : (-27'h8)) * (w3 & (25'h15))), (26'h1d), w4, (~^$unsigned((-9'h16))), {(5'h3), w7, (7'h1a), (-22'h18), w5, (10'h12), w8, (-30'h19), w10, (28'h15), (10'h17), (2'h3), (23'h12), (11'h15), w95, w1, (24'h15), w2, (26'h1), w95, w1, w98, w1, w7, (-6'h9), w99}, {(5'h1d), (20'h13), (-27'h1d), (-26'he), (17'he), w5, (-30'h2), w96, (6'ha), (2'h19), w7, (8'h1), w2, w4, (1'h1), (3'h15), w9, w9, (11'he), (-4'ha), (3'h6), w4, (-21'h11), w1, (3'h8), (29'h7), (-3'h11)}, (((-30'h8) <= (-14'h8)) ? (w8 ? (22'h18) : w5) : (-18'h3)), ((w3 << (-25'h15)) ^~ (w8 <<< w96)), w5, (-1'h10), $signed((~|(22'h4))), {w1, w7, w4, (24'h1a), (-22'h9), (23'h5), (-8'h6), w1, (-6'h19), (-3'hf), (-22'h0), (15'h1a), (-26'hf), (-19'hf), w96, (29'h1b), w8, (15'hb), (28'h14), (-22'h18), w3}, $unsigned(((12'h1b) << (26'ha))), $unsigned(((-8'h1e) >> w8)), (^(~|w8)), $signed((10'h16)), w9};
assign w95 = w9;
assign w96 = $signed((|($signed(w5) ? (-24'h7) : ((15'h8) <<< {(-23'h1b), (19'he), w1, w5, w9, (6'h13), (2'h9), (-23'h9), w5, w9, (6'h17), w6, (-8'h0), w5, (-2'h2), w6, w1, (17'h1a), w100, w100}))));
assign w97 = ({$unsigned(w98), (~&(14'h2)), $signed(w3), ((12'h7) >> w2), (^w10), $unsigned(w99), (w8 && (-25'h1)), {w99, (-27'h11), (-8'h1d), w7, w1, (-25'h17), w6, (26'h1b), (-15'h11), w9, (-2'h7), (-26'h14), (27'h17), (9'h17), w100, (3'h3), w9, w6, w98, (-22'h18), (15'he), w1, (1'hf)}, {w5, (-9'h4), w3, (-29'h18), w5, (-1'h1a), w9, (-8'h14), w98, (-9'hb), (19'h2)}} ? w5 : $unsigned($unsigned(w8)));
assign w98 = (~&{((22'h5) ? w4 : w3)});
assign w99 = ($signed((~|{w2, (-21'h15), (23'hc), (31'h1a), w4, w8, (-9'h1a), (-22'he), (24'h5), w10, (10'h13)})) <<< (^(w100 == (w10 ? w4 : ((-9'hb) ? w4 : (15'h14))))));
assign w100 = ({w10, $unsigned((-5'h8)), (w6 ? w8 : (1'h8)), ((-5'h1e) ? (-6'h13) : (-2'h1b)), $signed((-16'h16)), w2, (~|w1), {(5'h13), (-13'hd), (-9'h15), w4, (-9'h14), w7, (17'h5), (-27'h1c), w8, w4, w3, w6, (17'hb), (30'ha), (-10'h8), (11'hd), w10, w6, w4, (-13'h5), w10, (-25'h11), (-16'h11), w5, (27'h5)}, ((30'hd) ^~ (-21'hc)), $signed(w3), ((30'h1a) <= w4), {w2, w4}, (-4'h1), (w3 * (-15'h1a)), (w2 ? (-3'ha) : w10), {w5, w7, w2, w6, w6, (-18'h18), (-4'h1a), (-5'hc), (-2'h0), w5, w2, (28'he), (3'hc), w7, (34'h1a), (-14'h10), w1, w9, (-7'h6), (20'hb), (-31'h1c), (4'h9), w9, w3, (23'hb), w6, (-31'h1a)}, {(-21'h1c), (-30'hc), (28'hc), (20'h18), w4, (-23'h14), (19'h7), w4}, (27'hb), w8} ? ((^((-1'h9) ? w8 : w5)) ^~ (!$unsigned($unsigned((24'ha))))) : $signed((-(((29'h9) > (-3'h3)) === {w5, w8, (-28'h10), w2, (23'h11), w4}))));
assign y = {w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100};
endmodule
