module test_module(y, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10);
output wire [1458:0] y;
input wire [26:0] w1;
input wire [24:0] w2;
input wire [23:0] w3;
input wire [1:0] w4;
input wire [5:0] w5;
input wire [12:0] w6;
input wire [27:0] w7;
input wire [16:0] w8;
input wire [14:0] w9;
input wire [13:0] w10;
wire [10:0] w11;
wire [2:0] w12;
wire [11:0] w13;
wire [6:0] w14;
wire [14:0] w15;
wire [9:0] w16;
wire [9:0] w17;
wire [10:0] w18;
wire [25:0] w19;
wire [4:0] w20;
wire [27:0] w21;
wire [2:0] w22;
wire [14:0] w23;
wire [11:0] w24;
wire [8:0] w25;
wire [29:0] w26;
wire [14:0] w27;
wire [8:0] w28;
wire [25:0] w29;
wire [15:0] w30;
wire [16:0] w31;
wire [1:0] w32;
wire [18:0] w33;
wire [25:0] w34;
wire [17:0] w35;
wire [20:0] w36;
wire [25:0] w37;
wire [6:0] w38;
wire [7:0] w39;
wire [4:0] w40;
wire [22:0] w41;
wire [20:0] w42;
wire [8:0] w43;
wire [29:0] w44;
wire [5:0] w45;
wire [25:0] w46;
wire [15:0] w47;
wire [11:0] w48;
wire [11:0] w49;
wire [4:0] w50;
wire [21:0] w51;
wire [5:0] w52;
wire [6:0] w53;
wire [25:0] w54;
wire [15:0] w55;
wire [26:0] w56;
wire [27:0] w57;
wire [27:0] w58;
wire [25:0] w59;
wire [4:0] w60;
wire [1:0] w61;
wire [23:0] w62;
wire [29:0] w63;
wire [17:0] w64;
wire [13:0] w65;
wire [25:0] w66;
wire [13:0] w67;
wire [20:0] w68;
wire [4:0] w69;
wire [24:0] w70;
wire [16:0] w71;
wire [26:0] w72;
wire [23:0] w73;
wire [1:0] w74;
wire [25:0] w75;
wire [25:0] w76;
wire [10:0] w77;
wire [7:0] w78;
wire [25:0] w79;
wire [15:0] w80;
wire [19:0] w81;
wire [28:0] w82;
wire [22:0] w83;
wire [11:0] w84;
wire [3:0] w85;
wire [8:0] w86;
wire [17:0] w87;
wire [4:0] w88;
wire [10:0] w89;
wire [22:0] w90;
wire [21:0] w91;
wire w92;
wire [21:0] w93;
wire [17:0] w94;
wire [25:0] w95;
wire [23:0] w96;
wire [12:0] w97;
wire [10:0] w98;
wire [24:0] w99;
wire [7:0] w100;
assign w11 = w65;
assign w12 = (!((|{(4'h17), (10'h9), w27, w19, w82, w100, (-12'h1d), w85, w99, w22, w76, (-4'h0), w53, (2'hc)}) ? w16 : $unsigned(((w7 ? w42 : w93) ^~ (^~(3'h1b))))));
assign w13 = $signed({(w63 != (-15'h6)), (17'h1), ((19'h1b) ? (28'h14) : w4), (^w6), (-10'h16), ((17'h1) <<< (8'h15)), (w99 ? w16 : w46), (+(6'ha)), (w44 >= w20), (w58 !== w53), ((10'h6) !== w62), (w26 != (29'h1e)), $signed(w74), {(20'h12), (6'h10), (-26'h3), (13'h15), (4'h1c), (-26'h7), w74, w95, w62, w21, w73, w1, w93, w83, (-15'h16), w59, (-29'h1), w61}, ((10'h15) || (-19'h1c)), (w82 ? w15 : (-24'h10)), (+w97), (18'h2), ((1'he) ? w52 : (-4'h1a)), (w38 ? w92 : w57), {w100, (-6'h3), w100, w19, (-31'h16), (30'ha), w55, (-22'h18), w49, (22'h8), w67, w19, (2'h10), (-25'h7), w60, w79, (15'h6), w24, (17'h18), (-29'hd), w65, (-29'h16), (5'h1c), w32, (-6'h14), w91, (-28'hd)}, {(-27'h4), (8'hc), w30, w67, (3'h13), w27, (9'h3), w57, w44, w53, (1'hd), w93, w85}, w4, {(11'h2), w95, w83, (9'h8), (30'h2), w3, w66, w68, (-10'h1b), w80, (5'h16), (-5'h1), (24'h2), (25'h16), (27'h11), w47}, ((-10'h15) >> (-9'h8))});
assign w14 = {{(-25'h6), w22, w82}, w49, {(-9'h0), (19'h1), (-24'h7), w41, w43, w24, w46, w91, w76, (20'h7), (-23'h14), w43, w87, (-27'h10), (30'h2), w87, w79, w43, (-28'h0), w23, (-30'h18), w7, w63, (-20'hd), (18'ha), w55, (19'h10)}, (-w69), (w59 ? (19'h1b) : (w35 ? (22'h1c) : (-13'h1))), ((|(12'h8)) ? ((30'ha) ? w56 : (23'h1c)) : (15'h19)), $unsigned($signed(w75)), (30'ha), (^~$unsigned(w50)), {(-23'h13), w88, w52, w53, w84, w79, w78, w4, w79, w31, w82}, w78, w72, $signed((-23'h5)), $unsigned((&w88)), (-22'h18), (24'h15), (^((-19'h9) ? (9'h19) : w42)), $signed($signed(w36)), (-22'h1), (((16'he) ? w85 : w42) ? (w2 & w6) : (|(30'he))), (-25'hc), w84, ((-30'h0) ? (w67 && (-18'h2)) : (w33 & (11'h15))), ((-27'h1) ? (~&(6'h19)) : (12'h19))};
assign w15 = $unsigned(((+((-7'h2) >= w62)) ? (-27'hd) : (w37 ? (6'h1d) : (-13'h1c))));
assign w16 = ((~^(((19'h1d) ? w97 : (-9'h2)) >= w80)) ? {(-21'h13), $signed(w18), w28, (w17 ? w89 : w23), (|(-19'h6)), (w44 * (-25'hc)), w76, (w63 <= (-18'h1b)), {w29, (2'h4), w60, w55, w58, (26'h1e), (-2'h0), (-11'hd), (-7'h1a), w85, w59}, {(9'h10), w31, w35, (-8'he), w35, w36, w68, (-30'h2), w49, w89, w90, w3}, (w19 > (-10'h2)), {(-11'h16)}, (-w94), w80, {(-9'h13), w71, (1'h1a), (5'h1b), w38, w9, (25'h19), (7'h1), w67, (31'h17), w5, w74, (-16'h17), (31'h1c), (12'h1c), (-23'h19)}, {w60, w18, w57, w7, w64, (8'h1a), (1'h10), (-32'h3), (-23'h1b), (-19'h1a), (-1'h3), w48, w51, w54, (-10'h19)}, (|w29), (+(12'h1a)), (w94 ? (-26'h15) : w39), (!(5'h11)), {w22, w8, w29, (-16'hf), w18, w87, (7'h3), w63, w30, w59, w40, w37, w6, (-18'h1), w60, w39, w90, w7, (-26'h16), (2'h6)}, $unsigned((26'h10)), (-19'he), (|w97)} : {((6'h12) ? w52 : (-9'h4)), (+w70), w56});
assign w17 = ({(-39'h7), {w77, w81, w24, w47, w4, (30'h12), w20, (12'h3), (10'hf), w56, w64, (8'h1d), (-3'hf), (17'h1), w28, w83, w95, w9, (18'h1e), (-4'h1a)}, (23'h1e), $signed(w42), $signed(w60), (~^w31), $signed((-22'h8)), ((13'h17) >= w57), ((-22'h9) >>> (6'h7)), w68, (|w62), ((-30'h19) ? (2'h5) : (-11'h1c)), (-19'h16), $signed(w61), ((15'h7) && w80), $signed(w1), {w29, (2'h1c), w39, w23}, (~&w38), w18, $unsigned(w73), ((-20'h5) ? w61 : (-30'h9)), (w65 && (-22'h3)), (+w31), ((30'h1c) ? (28'h4) : (-10'h1d)), (w55 && (21'hd))} ? $unsigned($unsigned($signed((w97 | (-3'h8))))) : (~^(25'ha)));
assign w18 = ({$signed(w65), (w70 ~^ (-7'h7)), (w76 ? w86 : (-6'h8)), ((23'h3) ? w28 : (3'h11)), (-12'h1c), (&w49), $signed(w90), ((32'h6) ? (-26'h5) : (14'h6)), (-14'h18), (17'h14), {w82, w31, w29, (9'hb), (-15'hd), (17'h1d), (-13'hb), w71, w65, (16'h1d), w32, w37}, $signed((-13'h13)), ((-5'h1e) * (13'h1e)), $unsigned((6'h1b)), (~^(-4'h13)), $unsigned((-4'h11)), {w94, w99, w78, (1'h1d), (16'h9), w4}, w81, (19'h1d), w80, (-29'h18), ((-16'he) >> w56)} ? (-6'h10) : (4'h1e));
assign w19 = w21;
assign w20 = (~^(+w36));
assign w21 = w61;
assign w22 = w2;
assign w23 = (~|(18'h1));
assign w24 = (-(14'h13));
assign w25 = ($signed((19'h11)) ? (17'h17) : (^~(~&$unsigned((-2'h10)))));
assign w26 = ({(w71 ? (3'h17) : (-11'h8)), w90, w91, (~^(5'h12)), {(11'h8), (-16'hf), w46, w77, w1, (-17'ha), (27'h15), w37, w34, w73, (1'h15), (24'hc), w56}, (2'h3), ((-16'h19) ? w77 : w7), {(-9'h6), (3'hb), (24'h11), (-28'h2), w63, (8'h13), w33, w43, w93, w99, w58, (13'he), w86, (-7'h16), w83, (18'h18), (-28'h5), (22'h1e), w47, w81, (-17'h1c), (16'h16), (-24'h1d), (4'h1e), (-16'h10), w57, (7'h19)}, (18'hb), w35, {w95, w76, (10'h18), (-3'h5), (7'h14), w74, w61, (-25'h1d), w100, w46, (-23'h18), w81, w2, w89, w81, w47, w64, w100, (-21'hf), w10, (26'hc), w82, (13'h8), (8'h12)}, {(-1'h3), (26'h6), w28, w63, (9'hd), (-22'h2), w2, (10'h17), w77, (-4'h18), w39, w64, w29, (-28'hd), w27, (18'h9), w60, (15'h1), (-10'h9)}, (w33 + w55), (-29'h7), w27, (w28 ? w32 : w47), {w49, (27'hc), w78, (-9'h11), w4, (-8'h17), (-24'h18), (-7'h6), w100}, (23'hd), (27'h11), w64, w96, $unsigned(w93), w76, (~|(-21'h9))} == (w7 ? $signed((w45 * $unsigned(w61))) : $signed((~^$signed((9'h17))))));
assign w27 = w58;
assign w28 = {((-7'h1d) ^~ (!(5'h5))), ((-22'h1c) ? (10'h1c) : {(17'h1b), (8'h1), (30'h15), w61, w53, w68, w68, (6'h14), w33, (19'h12), w95, (28'h3), (15'h7), (5'h1a), w38, (-27'h5), w88, (-17'hb), (24'h1e), w51, (-3'he), w52, (6'hb), w65, w49, (-3'h18)})};
assign w29 = ({(w93 ^ w53), (+w87), (-23'ha), (5'h5), {(-27'h11), (15'h2), w4, (-18'h10), (10'h11), w98, w96, w83}, (w32 ? w84 : (-23'h16)), (^w41), ((-6'h1e) || w68), (-17'h1), $unsigned((-3'h1b)), (w54 ? w80 : (29'h1)), (w83 ? w89 : w84), w46, $signed(w99), $unsigned(w72), (+w67)} << $signed((~&(-26'h2))));
assign w30 = $unsigned((((^(10'h1c)) ^~ {(9'h1d), w86, (26'h7), (26'h7), w38, w91, w41, (6'ha), (-8'h1d), w83, (-8'h8), w64, w9, w33, w37, (22'h14), (8'h14), (7'hb), w78, w8, (-20'h2), w33, (-14'h1), w77, (22'hb), (13'h1d), w81, (-25'h1e), (-19'h18), (-19'h1e)}) ? (((4'h1) ? w38 : (5'h14)) >>> $unsigned((&(24'he)))) : $unsigned((+(w73 ? (-8'hb) : (-30'he))))));
assign w31 = (w41 !== (~^({(27'h1a), w84, w68, w46, w45, (9'h14), w97, (-13'h16), (4'hf), (-15'h15), (9'hf), w3, w89, (22'h1), (-9'h10), (6'h17), (-29'h18), (29'hd), (15'h2), w47, (3'h5), w48, (2'h1a), w55, (30'h4)} >> ($unsigned(w33) ? (!(27'hd)) : (~^(24'h1a))))));
assign w32 = (11'h9);
assign w33 = (((~^{(-19'h19), w66, (-8'h7), w6, (15'h11), w67, w66, w37, (-10'hc), w99, w80, (-23'h13), (14'h6), w55, w5, (-22'h13), w98, w2, (22'h10), (17'h12), w62, w44, (3'h12)}) || {(-9'h5), w40, (7'h1e), (27'h17), (-10'hc), w66, (-1'h1c)}) === ($signed((((20'h1) ? (-28'h1a) : (-31'h12)) << (^~(-7'h4)))) ^ ((-23'h8) + w98)));
assign w34 = ({(~|w5), $unsigned(w58), (w3 ? w67 : w55), (!w67), ((-22'h17) == w7), $unsigned((-5'hd)), (3'h8), w81, $signed((20'h17)), $signed(w45), w66, (w74 ? (10'h8) : w49), {w5, w51, w84, (13'he), (24'h7), w1, w65, (18'h2), w95, w72, w10, w95, w92, w1, (3'h13)}, (5'h15), (w84 ? w6 : (26'h16)), w66, ((-6'h1d) ^~ w47)} ? ((21'h8) === (-5'h5)) : $unsigned($unsigned({w75, w72, (-30'h0), (24'ha), w84, w89, w6, (-2'h12), w37, w1})));
assign w35 = w44;
assign w36 = ({{w4, w52, w5, w51, (-31'h2), w54, (18'hb), (-2'hc), w75, (25'h1), (18'h1e), (-4'h1), (-25'hb)}, w46, (w96 ? w59 : w80), ((-11'h16) - (30'hb)), w79, w88, w81, w46, (-13'h1e), (w66 + w3)} || ($signed((((-22'hf) !== w99) ? (w59 ? w67 : (-5'h2)) : (!(15'h1a)))) > ({(2'h17), (-14'hf), w39, w70, w75, (29'h16), (12'h18), w74, w94, (-21'hb), w6, w95, (-14'h10)} <<< (((-1'h9) ? (-15'h12) : w10) ? ((-22'h1b) ? w54 : w81) : (w38 ? w86 : (8'h1))))));
assign w37 = $unsigned((~&(-8'h1e)));
assign w38 = (^(({w41, w69, w7, w6, (15'hf), w63, w43, w6, w57, w68, (-5'h6), (8'hc), (26'h4), (-29'h9), (-11'h13), w53, w56, w47, w98, (-31'h19), (-14'h9), w10, w92, (13'h3)} ? (~&w89) : $signed(w61)) ? (-1'ha) : (2'h1e)));
assign w39 = w66;
assign w40 = $unsigned({((22'h13) ? (-5'h1c) : w81), {(28'h14)}, (w8 ? (33'h4) : w75), $signed((-21'h13)), (-19'h1e), $unsigned((-21'ha)), (~^(3'h16)), (w95 != (12'h1a)), ((23'h6) ? (-25'h11) : (15'h1a)), w42});
assign w41 = ({$unsigned(w42), (9'ha), {(-10'h2), w45, w7, (-3'h12), (15'hc), (-24'h19), (6'h17), (31'h8), w66, (14'hc), (11'h5), (-20'ha), w79, (-23'h1e), w7, w80, (8'h18), w92, (-30'h1a), w1, (-29'h1d), (7'h19), (30'h2), (23'h15), w43, (23'h1b), w51, (30'h12)}, ((-11'h17) >> (27'h19)), (w61 ? w87 : (13'he)), (^~(-24'h1a)), $unsigned(w56), (w60 + w76), ((-28'h10) ? (-19'h16) : (-20'h6)), {w51, w56, (-17'hb), (-28'hf), (25'hb), (-18'h8), w73, w83, (25'h1a), (9'h3), (25'hd), (-31'hb), (19'ha), (-5'h5)}, $signed(w45), (~^w86), ((-17'hf) ^~ (-7'h1)), (w56 ? (-21'h18) : w72), (w91 ~^ (4'h4)), (&(-22'h4)), (w84 === (1'h4)), (15'hd), ((16'hb) | (2'h5)), w71, $unsigned((-14'h1d)), $signed((25'h18)), {w54, w52, (17'h1c), w89, (-12'ha), (-8'h0)}, $unsigned((10'h6)), {w72, w98, (11'h7), w65, (12'h1b), (-19'hb), w55, w87, w5, (2'h1e), (-3'h4), w79, (-24'ha), (6'h10), (2'h5), (12'h1e), (21'h4), w3, w53, (-6'h1b), (-28'hb), w5, w68, (11'he), w77, w76, w67}} ? (((13'h19) || {w59, w2, w53, w44, (-13'h12), w65, w88, (25'h1), w82, (-29'ha), (-27'h3), w83, (15'h1a), w3, (-4'h4), w98, (-29'ha), w75, w45, w42, (-11'hf), (-26'hb), w97, w82, (-24'h1a), (24'h4), (8'hc), w60}) ? w53 : {w77, (-28'h1c), (-23'h11), w8, w43, w89, w64, w65, (20'h18), w96, w50, w49, w50, (1'h14), w44, (24'h1c), w55, w58, w87, (-12'h12), (18'h16), w62, w56, (21'h12), w99, w4, w59, w70}) : $signed((+{(26'h1a), w99, (-9'h17), w75, w5, (-26'h1), (2'h13), (29'h12), (21'h15), (-8'h1c), w48, w49})));
assign w42 = (^(22'h7));
assign w43 = $unsigned(w81);
assign w44 = w46;
assign w45 = ({$signed((-26'hc)), (-17'hd), (-(-3'h12))} ? ({(24'h13), w96, (-9'h11), (-21'h1b), (-29'hc), (6'hc), (-29'h11), (22'hc), w61, w68, w10, (-3'h17), w93, (-21'hf), (6'h5)} >>> ((-5'h4) || (~^(-(-19'h1e))))) : (~^(((1'hd) ? w59 : (19'hd)) << (w67 ? w60 : w90))));
assign w46 = ((-(({(-24'h17), w94, w97, (-28'hb), w85, w50, w92, w70, w74, (25'h7), (-25'h2), (-25'h5), w62, (-9'hc), w87, (28'hd), (-16'h4), w100, (-29'h5), (31'h2)} > (w55 << w56)) ? w49 : (w61 ^ {(-15'h16), (-6'h8), w62, w78, (-12'h0), w100, (-23'hc), w90, (19'h17)}))) <<< (-9'h12));
assign w47 = (~&(($unsigned((-33'h10)) ? (15'h1c) : $signed((-7'ha))) ? {w52, w75, (28'hb), w75, w62, w70, (13'h4), (19'hc), (-30'h0), w50, (-16'h1d), (8'h13), (-15'h8), w90, w90, w62, (28'h10), (-3'h13), w4} : {w72, (-20'hb), w81, (-32'h16), (10'ha), w70, w68, w98, (1'h3), (14'hf), (-21'hc), w62}));
assign w48 = (^~(($signed((+(-27'h17))) >>> (~&(31'h13))) ? ((^(22'hd)) >>> $unsigned((w65 ? (26'h1a) : w10))) : (w50 ? {(-22'h1a), w64, (28'h12), w82, (-28'h3), w64, w54, (-19'hf), (-1'hc), (-18'h11), (26'h1b), w97, w56, (-24'h1a), (20'hf), w57, (23'h9), (-4'h19), (-31'h1d), w7, w4, w96, w78, (22'h1c), w96, w58, (-14'h19), (-13'h1a), (16'h1e)} : (+(17'h5)))));
assign w49 = w58;
assign w50 = ($unsigned($unsigned(({w57, w70, (-2'h19), w78, (2'h1d), (-13'h12)} ? {w73, (-6'ha), w63, w53, w51, w72, (13'h3), w75, w65, w68, (-18'h6), (-30'h0), w63, w99, w90, w75, w62, (-8'h16), w93, (-26'hf), w82, (-23'h1d), w61, w80, w8, (-7'h10)} : (|(-29'h14))))) - $unsigned((&((w4 ? w91 : (6'h1a)) >> ((4'h15) ? (-8'he) : w67)))));
assign w51 = (24'h7);
assign w52 = (w8 >>> {((-7'h15) < (4'hf)), (w96 === (-28'h18)), (20'h18), (^w77), $unsigned((-28'hb)), (|w84), (7'h1), w56, (-8'h16), (w1 >>> (-1'h1)), (w73 ? w76 : w56), w88, (^~(19'h17)), {w87, w82, (-4'h11), w63, (6'h14)}, w1, w79, (^w63), (w62 ? w76 : w98), ((30'h1d) ? (20'h1d) : w62), w53, $unsigned((26'h1a))});
assign w53 = {w93, w54};
assign w54 = w60;
assign w55 = ({w66, ((28'hb) ? w59 : w59), {(28'h1a), w66, w63, w68, w72, w70, w99, (23'h11), w4, (-2'he), (-26'h2), w1, w84, (12'h5), w5, w100, (8'h13), (-9'h12), (7'h4), (-22'h1c), w64, (-25'h1)}, ((5'h18) === w67), w61, ((-9'h14) ? w56 : w98), {(7'h14), w73, (-13'h9), w100, (-12'h1c), (26'h3), w61, w79, (-32'h6), (-24'he), w62, w69, (-30'h19), (-17'hc), w90, (-18'hf), w85, (-24'h19), w77}, (22'h1d), w96, (+w57), (~^(8'h8)), (|(9'h5)), (14'h6), {(-3'h3), w92, (1'h14), (20'h3), (8'h3), w65, w76, w95, w8, w76, w100, (-18'h1e), w70, (12'ha), w1}} || {w97, $signed(w64), w71, (5'h7), w6, w56, (w77 ? (16'he) : (28'ha)), (16'h12), (|(19'h1c)), $signed(w70), (^(-6'h8)), ((8'h15) ? w72 : (-5'h10)), {(-16'h4), (-4'h1d), (18'h19), (10'hf), w91, (-19'h10), w99, w97, w90, (27'h1e), (21'ha), w81, (26'h6), w75, (19'h1b), w79, w74, (-14'h1), w73, w96, w77, w62, w68, w97, (-23'h18), w60}, ((-21'h15) <= (18'he)), {(-32'hf), w81, w60, (4'h15), (28'h7), w62, w76, w71, (8'hc), w100, (-19'he), (22'hc)}, (+(-3'h13)), ((-6'h1b) ? w61 : w77), {(-13'h10), w89, (23'h1d), (-25'h9), w92, w88, w57, w97, w3, (8'hb), w80, (11'hb), (-26'hd), (-15'h9), w10, w56, (-16'ha), w58, (28'h1b), (7'h1a)}, $signed((12'h4)), (-17'he), (w8 ? w80 : (-15'h1d)), (~|(16'h13)), ((29'hf) != (14'h5)), $signed(w9), (-21'hc), (-9'h17), $signed(w70)});
assign w56 = $signed((-22'h0));
assign w57 = ((-31'h0) ? (3'h8) : (({(29'h19), w98, w63, w71, (-17'h4), (-4'h12), (18'h11), w58, (7'h13)} >> ((6'hf) && w61)) ? w58 : (-28'h10)));
assign w58 = (~&(-3'h16));
assign w59 = ({$unsigned(w68), (w99 >= w9), w80, (-17'h5), $unsigned((5'h8)), ((14'hb) ^ (28'h11)), $signed(w78), $unsigned(w84), $signed(w70), {(-28'hc), w71}, (~^w4), $signed(w86), (w89 === (-2'hc)), ((-28'he) >>> (1'h4)), w64, w97, (w99 >>> w79), (-1'h1b), ((28'hc) ? (-23'h3) : (-22'h12)), {(22'hc), (-22'h0), (-3'h7), (24'ha), (14'h1), (-2'h8), w63, (-16'h13), (-5'h12), w85, (-5'h10), w92, (17'h1e), w7, (21'h9), w62, w93, w69, w60, w94}, ((-30'h1) || w73), w86, ((32'hb) ? w62 : (-24'h10)), ((-19'hc) !== (10'h10))} >= w74);
assign w60 = ((~^(!$signed($signed(w95)))) | ((w95 === ($signed(w63) != w100)) !== (-7'he)));
assign w61 = w79;
assign w62 = $unsigned($unsigned(((-11'h12) ? w73 : ((w84 ~^ (8'h17)) <<< (~&w63)))));
assign w63 = (($unsigned((4'h14)) ? $unsigned((|(w70 !== (-19'h8)))) : w84) !== ({w79, (29'h4), w99, (9'h6), w81, (30'hc), (5'h1d), (6'h1), (-22'h2), w67, w69, w70, (5'h9), w9, (-32'h7), (15'h14), w6, w83, (29'h9), w70, w96, (30'h2), w4, w67, w85, w99} >= ((^~{(-5'h6), (11'h1), w97, (-1'h9), w84, w65, (31'h8), (-10'h12), w5}) ~^ $signed((!w72)))));
assign w64 = (({w69, (17'h1c), w93, (3'h13), (25'h3), (25'h6), w67, w73, (22'he), w82, w68, w89, (-27'hb), (22'h2), w68, (-11'h17), (11'h17), (-26'h12), w100, w7, w83, w87, w96, (17'h13)} < (-{w91, (20'h8), (-4'h13), w70, (4'h15), (3'h17), w95, (7'h1d), w91, (18'h10), (-22'h5), w81, (-21'hd), (-23'h1b), w3, w66, w83, w84, w5, w79, w10, w4, (-29'hb), w79, (24'h17), w77, (26'h1), w77, w7})) ? (18'h14) : ((|$signed((-27'he))) ? $signed($unsigned(w6)) : $signed(((-3'h4) !== (-9'hc)))));
assign w65 = (({(-23'h0), w81, (13'h3), w88, w7, (29'h1e), w97, (7'h2), (-25'h1), (4'h7), w89, w69, (-6'he), (-22'h4), w7} != (&((~&w71) ? (+(-19'h1e)) : $unsigned((-22'hd))))) < $signed(((w3 ? w76 : (30'h14)) ? (~^w1) : ((28'h1e) ? w75 : w94))));
assign w66 = (~^(^~(5'h2)));
assign w67 = $unsigned($unsigned((~^{(-25'h3), w93, w86, (-7'h18), w1, (-4'h2), (-30'h6), (14'hb), w91, (15'h13), (22'h10), (-29'h1e)})));
assign w68 = w70;
assign w69 = ({((-1'h2) === w5), (w9 >> (7'hf)), (~|(6'h1)), ((21'h6) ^~ (13'h1)), (|w95), ((-4'h18) ? w99 : (-16'hb)), {w71, w93, w81, (-11'h3), w88, (-23'h17), (9'h6), w7, (-30'h0), w79, w91}, (~^(-27'hd)), (^(11'h14)), $unsigned(w71), (~^w4), {w5, (-19'h2), w97, (7'hc), (-19'h7), (-4'h1), w1, w5, w94, (-12'h3), w100}, (w77 >>> w95)} ? ((w80 != (^((-17'h9) ? (24'h18) : (2'h1a)))) > (1'h16)) : (($signed(w77) ? {(17'h1d), (29'h1c), w77, (12'h9), w98, w85, w3, w88, w92, w93, w86, w79, w6, (-13'h18), w83, w75, w100, w92, (8'hc), w96, (22'he), w94, (25'h3), (13'h15), (1'hb), (-12'h5), (8'h1c), w97} : (~|(-20'h9))) ^~ {(-10'he), w91, w95, w90, (-3'h8), (29'h7), (-1'h4), w93, w70, w3, w100, w82, (-1'h7), w7, w72, w75, w77, (-14'h1), (-17'h10), (1'h16)}));
assign w70 = (-(-(~&((w95 ? w76 : w81) && (^(3'h18))))));
assign w71 = {(^~((-4'hf) ? (-1'hd) : (-17'h8))), ({(11'h11), (31'ha), (-12'h1e), (8'h15), w1, (21'h8), w72, (15'h17), w81, w93, (19'h8), (21'h12), w72, w100, (24'h1c), w87, (-13'h1d)} >>> ((-15'he) < w94)), (-15'h6), (w79 + {w95, (-12'hb), w87, (19'h9), w80, (-11'hc), w97, (24'h17), w82, w8, w76, w2, (2'h9), w72, (12'h12), w6, w72, w88, w80, w90}), (-2'h1d), $unsigned(((11'hc) <= (-21'h19))), (+$unsigned(w88)), (-1'h19), $unsigned($unsigned((-20'h1))), (32'h3), ((w87 & w97) + {(11'h18), (-4'h5), (3'h7), (-9'hf), (-23'h2), (-17'h1e), w3, w85, w92, (-24'h12), w96, (-8'h1e), w1, w73, w82, w84, w8, (8'h7), w87, w100, w73, w1, w72}), w77, ((w86 ? (-1'h11) : (-5'hc)) ? {w78, (14'h1d)} : (10'h3))};
assign w72 = w87;
assign w73 = (+({w95, (20'h17), w83, (10'h5), w85, (20'h16), (19'hb), (18'h1d), w2, w99, (-34'hd), w75, w88, (29'h3), w91, w74, w89, (14'h9)} + (!$signed($signed(w98)))));
assign w74 = (($signed(w93) ? (|(-25'h1a)) : {w3, (-1'h18), w93, (-29'h11), (3'h9), (-31'h1c), w87, (14'hb), w98, w86, (6'h4), w2}) ~^ (-30'h1a));
assign w75 = ({(-16'h6), w81, (w8 !== (18'h16)), (~|w5), w81, (&(27'h4)), {w95, (8'h6), w3, w83, w6, w83, (6'h9)}, w84, {w10, w85, w77, (23'ha), w6, (-23'hd), w82, w1, w7, w79, w99, (-27'hf), w89, (-16'h1), w2, w83, (5'hb), w97, (-11'h1d), (-19'h9)}, {w78, (-17'h3), w2, w80, w10, w100, (-18'h19), (-11'hb), w92, (-22'h5), w98, (-18'h4), (6'h12), (-18'h17), w94, w92, w94, (31'h18), (13'h12), w82, (-6'h19), w90, (-7'hc), (-6'h6), (-26'h2), w90, (27'h1c), (7'h10), w82, w96}, (~|w6), $unsigned((9'hd)), ((1'h2) ? (17'h19) : w98), ((-27'h7) ~^ w96), ((10'h3) >= (-5'h16)), {w96, w79, (-3'h1a), w89, w9, (-21'h10), (8'hc), (3'h15), (-1'h3), (16'h13), (6'h1b), w9, (6'hb), w4, (11'h1b), (17'h5), (33'h14), (15'h17), (-24'h4), (8'h7), (-28'h0), (-6'h9), (-15'h2), w9, w6, (-30'h12), w81, (6'h14), w91, (-7'h1c)}, $signed((17'h10)), ((18'h12) ? (24'ha) : w10), (-24'hd)} - {{(-8'h1b), w99, w3, w97, (-29'h10), w99, (-16'h3), w90, w85, (1'h6), w93, (-1'h1c), (18'h13), (-10'h2), w96, w78, (-17'h8), (7'hc), (-30'h6), w79, (4'hc), (-30'h1a), w90, (18'h5), (30'h7), w8, w88, (2'h4), w5}, {(-10'h6), (-5'h1), (31'h1), (13'he), (-10'h15), (7'h18), w88, (-12'h7), w5, w94}, ((-2'h19) << w8), {(-22'h5), (9'h1a), (11'h1), w7, (-20'h1a), w78, (-22'h1d), w4, w91, w8, w83, w85, (-30'h7)}, {w10, w90, w2, (-14'h5), w97, w8, (-24'h5), w79, (-14'hf), (4'h1a), (33'h11), (-2'h8), w85, (-9'h18), w96, w97, (21'h15), (17'h15), (-14'h10), w76, (23'h11), (1'h8)}, (~&(-29'hf)), (w5 & (31'he)), ((-15'h5) ^ w94), {w89, (20'h10), (-3'h10), w3, (26'he)}, $unsigned(w99), (-30'h5)});
assign w76 = {(-w4), (-26'h3), (20'h3), ({(22'h1b), (27'hd), w6, w7, w80, (-26'he), w81, w92, (6'h7), w5, (-26'h18), w85, (6'h17), w2, w78, w81} >> ((-6'h19) ? w88 : (-11'h16))), w100, ($unsigned((8'h9)) !== (w80 ? w97 : (-17'h1a))), ((w86 * w100) <<< {w5, w10, (24'ha), w6, (-21'h9), w84}), (-14'h13), (w88 >>> (w98 ? w1 : (14'h1a))), ({(20'hf), (-26'hf), (-22'h18), w91, w93, (11'h4), (20'h15), w7, w1, w82, w77, (27'h9), (2'hd), (-21'h1e), w6, w80, (-21'h18), (-10'hf), w2, (-31'hd), w77} ? ((25'h13) ? w86 : w79) : {(8'h8), (-21'h2), (-7'h1c), w98, (-17'h18), (-12'h16), (-21'h17), (-26'h1d), (-13'h1d), w88, (-21'h16), (-17'ha), (-7'h1), w82, w97, w2, w4, w8, w9, w89, (29'h19), (-24'hd), (23'h1e), w82, w10, (-24'h1a), w94}), (-19'h15), {w4, (-23'h1a), w9}, w10, (-25'h1e), (10'h8), $unsigned(((-6'h4) != (-6'h4))), {w96, (12'hc), w93, w89, w83, (-16'h3), (-11'hc), (-32'hc), w94, (-31'h1e), (3'h12)}, w97, ((w10 ? w3 : w86) ? {(20'h12), w100, w77, (-12'hd), (-7'h7), (5'h1e), w80, (1'hb), w89, (33'h1)} : (-4'hf))};
assign w77 = (w88 != (w94 >= (&w88)));
assign w78 = $unsigned((12'hf));
assign w79 = (-7'h16);
assign w80 = (+($signed(($signed(w4) ? (-29'hd) : w9)) ^ (+({(-25'h1a), w3, w91, w5, (-29'h1), (-5'h11), (19'h17), w10, (17'h10), (11'h8), w89, w9, (13'h3), (-2'h6), w1, (-11'h1b), (-25'h1d), (-6'h17), (19'ha), w83, w88, w87, (14'h2), (-12'h1d)} - $signed((7'hc))))));
assign w81 = w7;
assign w82 = $signed((~^(27'h10)));
assign w83 = (!w90);
assign w84 = w5;
assign w85 = $unsigned((-18'hb));
assign w86 = {(14'h9), $signed((-24'h10)), $unsigned((w92 ? (25'h13) : (-21'hd))), {w89, (-30'h10), w98, (-13'h9), (18'h8), w10}, w90, w1};
assign w87 = {w88, (16'h1c), ($unsigned(w98) - w2), ($unsigned((-26'h0)) ? (w100 ? w88 : (-21'hb)) : (21'hf)), (w98 > $signed((25'h1b)))};
assign w88 = (-10'h16);
assign w89 = (w95 >= ((~&(&{(13'h7), (25'h19), (-27'h4), (24'h17), w10, w1})) >> (23'hf)));
assign w90 = ({(^w91), (w4 + (-7'h12)), (w2 ~^ w99), w98, (w97 ? (-25'h10) : (19'h19)), (w5 * w92), (!(-18'h19)), (12'h1a), (-32'h1c), $unsigned(w93), $unsigned(w98), (|(29'hf))} ^~ (-$unsigned({w99, (1'h14), (8'ha), (15'h8), (-1'hb), w7, (11'h1d), w91, (-7'h1c), (-29'h4), w98, w96, w6, w5, (-10'h5), w93, (-14'h18), (7'h1e), w8, (-1'h1b), (13'h15), (22'h8), (-21'h17), w2, (-3'h1b), (-23'h12)})));
assign w91 = (&{{(12'h4), w98, w9, (-27'h1b), w5, w7, w99, (-4'h1b), (-1'h18), (-19'h4), w9, (28'h2), w94, (-1'h1a), w8, (20'h3), (-13'h2), (7'h16), (28'h1e), (24'h1d), w6}, w2, $signed((6'h5)), $signed(w4), $signed(w8), (|w6), $signed((25'h1)), (-13'h5), $signed((31'h1b)), (w7 === w92), {w4, w100, (29'h18), w3, w98, (-14'hb), w93, (-17'h5), (24'hc), (-15'he), (19'h13), w5, w3, w94, w92, w10, (8'h5), (-31'h5), (-23'h10)}, $unsigned(w10), $unsigned(w93), (w99 ? (31'hd) : w7), ((30'he) > (-17'h15)), ((-1'h1e) == w98), {w97, (27'he), (21'h1), (23'hb), (-9'h2), w10}, ((4'h3) ? w3 : (31'hd)), $unsigned(w99), w8});
assign w92 = ((($unsigned((^w100)) ? (^~w98) : (((-11'h9) <<< w3) > w6)) >= {w8, (-20'h12), w94, (3'h1a), (-15'h2), (-3'h6), (-10'ha), (7'h5), w5, (9'hc), (27'h17), w95, w5, (12'h7), w95, (-22'h15), w10, (-11'h19), (1'h11), w2, (16'h13), (-16'he), w96, w3, w4, w6}) > ((-{w93, w100, (-6'h0), (-13'h12), w94, (26'h12), (17'h7), w100}) != w9));
assign w93 = {{w9, w3, w2, (-11'h0), (-7'h9), w10, (-19'h1e), (-12'h9), w6, w2, (-12'hf), w94}, ((~|w3) ^ {w95, (-6'h9), (12'h8)}), (^~(w9 + w94)), ((w6 || w97) + $signed(w95)), {(-19'hd), w10, (1'h12), (32'he), w96, w99, w7, w95, w2, w1, (4'he), (33'h17), w98, (30'h6), (-24'h17), w6, (24'h10)}, (-w7), (-(&(35'h6))), $signed($signed(w94)), $unsigned((|w1)), $unsigned((~^(21'h3))), w4, ((w6 ? w4 : w96) + $signed((-16'h1e))), (w4 ? $signed((-1'h13)) : (w98 ? w1 : w6)), w99, (-9'h1b), (|w94), $signed(w4), {w96, (7'h1), w95, w9, w96, (-15'h2), w96, w99, w1, w96, (-31'h1c), w95, w6, w5, (26'h1a), w10, w96, (9'h18), w98, (11'hd), (24'h7), (26'hd), (20'h17), (-11'h1c), w99, (-18'hd), w4, w100}, (-15'h1), (-24'h19), $signed(w4)};
assign w94 = (~^(-10'h9));
assign w95 = w99;
assign w96 = {((2'h1d) ? w8 : (10'h1)), (|w3), (~|(w100 ? w1 : w1)), (32'h4), ((w8 ? w8 : (-21'h4)) ? {(-11'hb), w3, (-28'h9), w100, (-28'h18), (26'h12), w10, (16'h16), w98, (6'h2), (19'h16), (-18'h17)} : ((5'h3) ~^ (-15'he))), ((w98 && (28'h1c)) ^~ (!w98)), $unsigned((-27'he)), (~^(30'h2)), (13'h1b), $signed((21'h13)), (&$unsigned((-23'h13))), {(-18'h10), (2'h10), (10'h1e), (-22'h10), w99, w8, (28'h1c), (26'he), w9, w100, (19'h1a), w1, (-19'h1c), (16'h2), (28'h3), w8, (-21'h15), w4, (31'h19), (4'h19), (7'he), (20'h16), (-22'h15), (2'he), w1, w1}, w97, $unsigned(w97), ({w100, w100, w8, (25'hb), (-12'h1c), (-13'h8), w97, (20'h12), w3, (-15'h15), w1, (-7'h0), w99, w4, w10, (12'h1b), w7, (17'hc), w10, (-27'h1c), w2, (-4'h5), w99, (-3'h13), (-14'h14), (-27'h8), w10} >= ((-30'hf) != w8)), (6'h1a), $unsigned((&w7)), $unsigned((^w100)), (23'h1d), (-29'h2), (((-24'ha) < w10) === (-28'h19)), w100, w6, $signed(w8), ((17'ha) ? (w8 ? w10 : (-8'h1c)) : (^~w6)), ({w100, (10'h12), (24'h19), w1, (20'h17), (18'h1d), (-7'hd), w99, w4, (-6'h1e), (21'he)} == (&(15'h18))), (-(-10'h1)), ({(6'hb), (-25'h3), w7, w10, w98, w2, w2, (17'h1c)} ? $signed(w6) : ((22'hd) | w10))};
assign w97 = $signed((8'h1b));
assign w98 = {((7'hd) ? ((7'he) ? w7 : w2) : (-12'h1e)), (24'h1), ($unsigned(w5) ? {w9, (13'h6), w1, (17'h5), (18'h1c), (12'h3), (11'h1c), w2, (1'h19), (30'hc), (9'h17), w100, w3, (-26'h6), w3, w8, w6, w5, (1'h3), w6} : (&(9'h2))), (w10 ? {(26'h9), (25'h1b), (6'hf), (3'h8), w1, (22'hb), w6, (21'h13), (15'h13), w1, w10, w10, (27'h6), (-8'h1d), w5, (33'h1), (-9'h1), (-7'h0)} : w1), ((w99 ? (-24'h1a) : (1'h19)) ? ((-4'h1e) ? (-13'h18) : (28'hc)) : w4), ((w4 + w8) ~^ $signed((-18'h1d))), (~^(-2'h0)), (w8 + w100), w9, ((-w2) <= $unsigned((26'h13))), $unsigned(w2), {w1, (19'h5), (22'h4), w5, w3, w5, w99, w6, (-12'h10), w8, (-27'h19), (-27'h1), w8, w7, w9, (-20'h9), w1, w4, (-29'h17), (-10'h1), (20'hb), (19'h11)}, {(28'h15), (-23'hb), (22'h1c)}, (~|w8), w99, w9, $signed({w6, (30'h6), w1, (13'h16), w4, (25'h8), w5, w7, w7, w8, (-24'h1e), (-12'h9), (-20'h4), w7, w2, w4}), ((w1 >= w1) < $signed((-1'h1))), (+$unsigned(w2)), w99, ({(-4'h14), (32'h1c), w2, w3, (-21'h5), (6'h13), (-24'h16), (-28'h10), (-14'hf), w9, (-21'hf), (-8'h7), (-10'h0), (-4'h13), (-8'h2), (-20'h1c), w99, w10, (-26'h5), w9, (15'hb), (-9'h1c), w6, (-6'h12), (-16'h5), (13'hf), w9, (-26'h16), (-20'he), (-5'h5)} ? (w7 && (-2'h7)) : (+w10)), w6, $unsigned((!w7)), w8, {(17'h16), w10, (-30'h18), w7, (8'h3), w99, (-13'h17), (-19'h1a), (-5'h14), (-29'he), w2}, ({w8, w8, w6, w2, (-6'h16), (-11'h17), (26'h1), (29'hc), (-12'h18), (7'h1), (-30'h0), (16'h1), w5, w5, w1, w100, w4, (-19'h1b), (-1'h19), (17'h2), (27'hf), (-20'h8), (20'h9), w10, w9, w8} ^~ $unsigned(w5)), (-11'h4)};
assign w99 = (!$signed((|{w7, w3, (11'h19), w4, w4, w10, (26'h13), (8'hb), (-27'h2), (-12'hf), w3, w2, (-30'he), w3, w7, w6})));
assign w100 = w8;
assign y = {w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100};
endmodule
