module test_module(y, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10);
output wire [1393:0] y;
input wire [8:0] w1;
input wire [25:0] w2;
input wire [24:0] w3;
input wire [16:0] w4;
input wire [29:0] w5;
input wire [28:0] w6;
input wire [21:0] w7;
input wire [22:0] w8;
input wire [29:0] w9;
input wire [20:0] w10;
wire [24:0] w99;
assign w99 = ({(17'h19), {w3, (5'h9), w4, (15'hc), (-(30'h18)), (-(5'h14)), (27'h15), (24'he), w10, w8, w2}, w4, w1, ((-(18'h13)) + (-(25'h9))), (~|w2), ((8'h1e) ? (-(17'hf)) : (-(13'h9))), (w7 <= (-(13'h6))), (-(23'hd)), (4'h13), (w8 >> (-(11'h14))), w3, w8, {(-(4'ha)), w8, w10, (21'h1e), (1'h0), w5, (-(18'h16)), (1'h0), (7'h6), (12'h5), (14'h13), (-(26'h7))}, (w6 ? w6 : (-(13'h13))), (w5 ? w10 : (1'h0)), w2, w4, (4'h5), (11'h15)} ? $signed((|(17'h1e))) : $unsigned((~^((-(7'he)) ^ {(1'h0), (-(7'h10)), (-(13'h7)), w9, w3, (-(10'h13)), (3'h17), w6, (21'h6), (-(29'h6)), (28'h19), w1, (-(19'hf)), w10, (7'h12), (26'h9), w7, w6, (1'h0), (-(21'h15)), (18'hb), (-(6'ha)), (16'h16), (12'h17), (-(6'h17)), (-(7'h15)), w1}))));
assign y = {w99};
endmodule
